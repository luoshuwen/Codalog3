% generate problem of size 10000
reachable(X,Y) :- edge(X,Y).
reachable(X,Y) :- edge(X,Z), reachable(Z,Y).
increasing(X,Y) :- edge(X,Y), lt(X,Y).
increasing(X,Y) :- edge(X,Z), lt(X,Z), increasing(Z,Y).
edge(0, 1).
edge(1, 2).
edge(2, 3).
edge(3, 4).
edge(4, 5).
edge(5, 6).
edge(6, 7).
edge(7, 8).
edge(8, 9).
edge(9, 10).
edge(10, 11).
edge(11, 12).
edge(12, 13).
edge(13, 14).
edge(14, 15).
edge(15, 16).
edge(16, 17).
edge(17, 18).
edge(18, 19).
edge(19, 20).
edge(20, 21).
edge(21, 22).
edge(22, 23).
edge(23, 24).
edge(24, 25).
edge(25, 26).
edge(26, 27).
edge(27, 28).
edge(28, 29).
edge(29, 30).
edge(30, 31).
edge(31, 32).
edge(32, 33).
edge(33, 34).
edge(34, 35).
edge(35, 36).
edge(36, 37).
edge(37, 38).
edge(38, 39).
edge(39, 40).
edge(40, 41).
edge(41, 42).
edge(42, 43).
edge(43, 44).
edge(44, 45).
edge(45, 46).
edge(46, 47).
edge(47, 48).
edge(48, 49).
edge(49, 50).
edge(50, 51).
edge(51, 52).
edge(52, 53).
edge(53, 54).
edge(54, 55).
edge(55, 56).
edge(56, 57).
edge(57, 58).
edge(58, 59).
edge(59, 60).
edge(60, 61).
edge(61, 62).
edge(62, 63).
edge(63, 64).
edge(64, 65).
edge(65, 66).
edge(66, 67).
edge(67, 68).
edge(68, 69).
edge(69, 70).
edge(70, 71).
edge(71, 72).
edge(72, 73).
edge(73, 74).
edge(74, 75).
edge(75, 76).
edge(76, 77).
edge(77, 78).
edge(78, 79).
edge(79, 80).
edge(80, 81).
edge(81, 82).
edge(82, 83).
edge(83, 84).
edge(84, 85).
edge(85, 86).
edge(86, 87).
edge(87, 88).
edge(88, 89).
edge(89, 90).
edge(90, 91).
edge(91, 92).
edge(92, 93).
edge(93, 94).
edge(94, 95).
edge(95, 96).
edge(96, 97).
edge(97, 98).
edge(98, 99).
edge(99, 100).
edge(100, 101).
edge(101, 102).
edge(102, 103).
edge(103, 104).
edge(104, 105).
edge(105, 106).
edge(106, 107).
edge(107, 108).
edge(108, 109).
edge(109, 110).
edge(110, 111).
edge(111, 112).
edge(112, 113).
edge(113, 114).
edge(114, 115).
edge(115, 116).
edge(116, 117).
edge(117, 118).
edge(118, 119).
edge(119, 120).
edge(120, 121).
edge(121, 122).
edge(122, 123).
edge(123, 124).
edge(124, 125).
edge(125, 126).
edge(126, 127).
edge(127, 128).
edge(128, 129).
edge(129, 130).
edge(130, 131).
edge(131, 132).
edge(132, 133).
edge(133, 134).
edge(134, 135).
edge(135, 136).
edge(136, 137).
edge(137, 138).
edge(138, 139).
edge(139, 140).
edge(140, 141).
edge(141, 142).
edge(142, 143).
edge(143, 144).
edge(144, 145).
edge(145, 146).
edge(146, 147).
edge(147, 148).
edge(148, 149).
edge(149, 150).
edge(150, 151).
edge(151, 152).
edge(152, 153).
edge(153, 154).
edge(154, 155).
edge(155, 156).
edge(156, 157).
edge(157, 158).
edge(158, 159).
edge(159, 160).
edge(160, 161).
edge(161, 162).
edge(162, 163).
edge(163, 164).
edge(164, 165).
edge(165, 166).
edge(166, 167).
edge(167, 168).
edge(168, 169).
edge(169, 170).
edge(170, 171).
edge(171, 172).
edge(172, 173).
edge(173, 174).
edge(174, 175).
edge(175, 176).
edge(176, 177).
edge(177, 178).
edge(178, 179).
edge(179, 180).
edge(180, 181).
edge(181, 182).
edge(182, 183).
edge(183, 184).
edge(184, 185).
edge(185, 186).
edge(186, 187).
edge(187, 188).
edge(188, 189).
edge(189, 190).
edge(190, 191).
edge(191, 192).
edge(192, 193).
edge(193, 194).
edge(194, 195).
edge(195, 196).
edge(196, 197).
edge(197, 198).
edge(198, 199).
edge(199, 200).
edge(200, 201).
edge(201, 202).
edge(202, 203).
edge(203, 204).
edge(204, 205).
edge(205, 206).
edge(206, 207).
edge(207, 208).
edge(208, 209).
edge(209, 210).
edge(210, 211).
edge(211, 212).
edge(212, 213).
edge(213, 214).
edge(214, 215).
edge(215, 216).
edge(216, 217).
edge(217, 218).
edge(218, 219).
edge(219, 220).
edge(220, 221).
edge(221, 222).
edge(222, 223).
edge(223, 224).
edge(224, 225).
edge(225, 226).
edge(226, 227).
edge(227, 228).
edge(228, 229).
edge(229, 230).
edge(230, 231).
edge(231, 232).
edge(232, 233).
edge(233, 234).
edge(234, 235).
edge(235, 236).
edge(236, 237).
edge(237, 238).
edge(238, 239).
edge(239, 240).
edge(240, 241).
edge(241, 242).
edge(242, 243).
edge(243, 244).
edge(244, 245).
edge(245, 246).
edge(246, 247).
edge(247, 248).
edge(248, 249).
edge(249, 250).
edge(250, 251).
edge(251, 252).
edge(252, 253).
edge(253, 254).
edge(254, 255).
edge(255, 256).
edge(256, 257).
edge(257, 258).
edge(258, 259).
edge(259, 260).
edge(260, 261).
edge(261, 262).
edge(262, 263).
edge(263, 264).
edge(264, 265).
edge(265, 266).
edge(266, 267).
edge(267, 268).
edge(268, 269).
edge(269, 270).
edge(270, 271).
edge(271, 272).
edge(272, 273).
edge(273, 274).
edge(274, 275).
edge(275, 276).
edge(276, 277).
edge(277, 278).
edge(278, 279).
edge(279, 280).
edge(280, 281).
edge(281, 282).
edge(282, 283).
edge(283, 284).
edge(284, 285).
edge(285, 286).
edge(286, 287).
edge(287, 288).
edge(288, 289).
edge(289, 290).
edge(290, 291).
edge(291, 292).
edge(292, 293).
edge(293, 294).
edge(294, 295).
edge(295, 296).
edge(296, 297).
edge(297, 298).
edge(298, 299).
edge(299, 300).
edge(300, 301).
edge(301, 302).
edge(302, 303).
edge(303, 304).
edge(304, 305).
edge(305, 306).
edge(306, 307).
edge(307, 308).
edge(308, 309).
edge(309, 310).
edge(310, 311).
edge(311, 312).
edge(312, 313).
edge(313, 314).
edge(314, 315).
edge(315, 316).
edge(316, 317).
edge(317, 318).
edge(318, 319).
edge(319, 320).
edge(320, 321).
edge(321, 322).
edge(322, 323).
edge(323, 324).
edge(324, 325).
edge(325, 326).
edge(326, 327).
edge(327, 328).
edge(328, 329).
edge(329, 330).
edge(330, 331).
edge(331, 332).
edge(332, 333).
edge(333, 334).
edge(334, 335).
edge(335, 336).
edge(336, 337).
edge(337, 338).
edge(338, 339).
edge(339, 340).
edge(340, 341).
edge(341, 342).
edge(342, 343).
edge(343, 344).
edge(344, 345).
edge(345, 346).
edge(346, 347).
edge(347, 348).
edge(348, 349).
edge(349, 350).
edge(350, 351).
edge(351, 352).
edge(352, 353).
edge(353, 354).
edge(354, 355).
edge(355, 356).
edge(356, 357).
edge(357, 358).
edge(358, 359).
edge(359, 360).
edge(360, 361).
edge(361, 362).
edge(362, 363).
edge(363, 364).
edge(364, 365).
edge(365, 366).
edge(366, 367).
edge(367, 368).
edge(368, 369).
edge(369, 370).
edge(370, 371).
edge(371, 372).
edge(372, 373).
edge(373, 374).
edge(374, 375).
edge(375, 376).
edge(376, 377).
edge(377, 378).
edge(378, 379).
edge(379, 380).
edge(380, 381).
edge(381, 382).
edge(382, 383).
edge(383, 384).
edge(384, 385).
edge(385, 386).
edge(386, 387).
edge(387, 388).
edge(388, 389).
edge(389, 390).
edge(390, 391).
edge(391, 392).
edge(392, 393).
edge(393, 394).
edge(394, 395).
edge(395, 396).
edge(396, 397).
edge(397, 398).
edge(398, 399).
edge(399, 400).
edge(400, 401).
edge(401, 402).
edge(402, 403).
edge(403, 404).
edge(404, 405).
edge(405, 406).
edge(406, 407).
edge(407, 408).
edge(408, 409).
edge(409, 410).
edge(410, 411).
edge(411, 412).
edge(412, 413).
edge(413, 414).
edge(414, 415).
edge(415, 416).
edge(416, 417).
edge(417, 418).
edge(418, 419).
edge(419, 420).
edge(420, 421).
edge(421, 422).
edge(422, 423).
edge(423, 424).
edge(424, 425).
edge(425, 426).
edge(426, 427).
edge(427, 428).
edge(428, 429).
edge(429, 430).
edge(430, 431).
edge(431, 432).
edge(432, 433).
edge(433, 434).
edge(434, 435).
edge(435, 436).
edge(436, 437).
edge(437, 438).
edge(438, 439).
edge(439, 440).
edge(440, 441).
edge(441, 442).
edge(442, 443).
edge(443, 444).
edge(444, 445).
edge(445, 446).
edge(446, 447).
edge(447, 448).
edge(448, 449).
edge(449, 450).
edge(450, 451).
edge(451, 452).
edge(452, 453).
edge(453, 454).
edge(454, 455).
edge(455, 456).
edge(456, 457).
edge(457, 458).
edge(458, 459).
edge(459, 460).
edge(460, 461).
edge(461, 462).
edge(462, 463).
edge(463, 464).
edge(464, 465).
edge(465, 466).
edge(466, 467).
edge(467, 468).
edge(468, 469).
edge(469, 470).
edge(470, 471).
edge(471, 472).
edge(472, 473).
edge(473, 474).
edge(474, 475).
edge(475, 476).
edge(476, 477).
edge(477, 478).
edge(478, 479).
edge(479, 480).
edge(480, 481).
edge(481, 482).
edge(482, 483).
edge(483, 484).
edge(484, 485).
edge(485, 486).
edge(486, 487).
edge(487, 488).
edge(488, 489).
edge(489, 490).
edge(490, 491).
edge(491, 492).
edge(492, 493).
edge(493, 494).
edge(494, 495).
edge(495, 496).
edge(496, 497).
edge(497, 498).
edge(498, 499).
edge(499, 500).
edge(500, 501).
edge(501, 502).
edge(502, 503).
edge(503, 504).
edge(504, 505).
edge(505, 506).
edge(506, 507).
edge(507, 508).
edge(508, 509).
edge(509, 510).
edge(510, 511).
edge(511, 512).
edge(512, 513).
edge(513, 514).
edge(514, 515).
edge(515, 516).
edge(516, 517).
edge(517, 518).
edge(518, 519).
edge(519, 520).
edge(520, 521).
edge(521, 522).
edge(522, 523).
edge(523, 524).
edge(524, 525).
edge(525, 526).
edge(526, 527).
edge(527, 528).
edge(528, 529).
edge(529, 530).
edge(530, 531).
edge(531, 532).
edge(532, 533).
edge(533, 534).
edge(534, 535).
edge(535, 536).
edge(536, 537).
edge(537, 538).
edge(538, 539).
edge(539, 540).
edge(540, 541).
edge(541, 542).
edge(542, 543).
edge(543, 544).
edge(544, 545).
edge(545, 546).
edge(546, 547).
edge(547, 548).
edge(548, 549).
edge(549, 550).
edge(550, 551).
edge(551, 552).
edge(552, 553).
edge(553, 554).
edge(554, 555).
edge(555, 556).
edge(556, 557).
edge(557, 558).
edge(558, 559).
edge(559, 560).
edge(560, 561).
edge(561, 562).
edge(562, 563).
edge(563, 564).
edge(564, 565).
edge(565, 566).
edge(566, 567).
edge(567, 568).
edge(568, 569).
edge(569, 570).
edge(570, 571).
edge(571, 572).
edge(572, 573).
edge(573, 574).
edge(574, 575).
edge(575, 576).
edge(576, 577).
edge(577, 578).
edge(578, 579).
edge(579, 580).
edge(580, 581).
edge(581, 582).
edge(582, 583).
edge(583, 584).
edge(584, 585).
edge(585, 586).
edge(586, 587).
edge(587, 588).
edge(588, 589).
edge(589, 590).
edge(590, 591).
edge(591, 592).
edge(592, 593).
edge(593, 594).
edge(594, 595).
edge(595, 596).
edge(596, 597).
edge(597, 598).
edge(598, 599).
edge(599, 600).
edge(600, 601).
edge(601, 602).
edge(602, 603).
edge(603, 604).
edge(604, 605).
edge(605, 606).
edge(606, 607).
edge(607, 608).
edge(608, 609).
edge(609, 610).
edge(610, 611).
edge(611, 612).
edge(612, 613).
edge(613, 614).
edge(614, 615).
edge(615, 616).
edge(616, 617).
edge(617, 618).
edge(618, 619).
edge(619, 620).
edge(620, 621).
edge(621, 622).
edge(622, 623).
edge(623, 624).
edge(624, 625).
edge(625, 626).
edge(626, 627).
edge(627, 628).
edge(628, 629).
edge(629, 630).
edge(630, 631).
edge(631, 632).
edge(632, 633).
edge(633, 634).
edge(634, 635).
edge(635, 636).
edge(636, 637).
edge(637, 638).
edge(638, 639).
edge(639, 640).
edge(640, 641).
edge(641, 642).
edge(642, 643).
edge(643, 644).
edge(644, 645).
edge(645, 646).
edge(646, 647).
edge(647, 648).
edge(648, 649).
edge(649, 650).
edge(650, 651).
edge(651, 652).
edge(652, 653).
edge(653, 654).
edge(654, 655).
edge(655, 656).
edge(656, 657).
edge(657, 658).
edge(658, 659).
edge(659, 660).
edge(660, 661).
edge(661, 662).
edge(662, 663).
edge(663, 664).
edge(664, 665).
edge(665, 666).
edge(666, 667).
edge(667, 668).
edge(668, 669).
edge(669, 670).
edge(670, 671).
edge(671, 672).
edge(672, 673).
edge(673, 674).
edge(674, 675).
edge(675, 676).
edge(676, 677).
edge(677, 678).
edge(678, 679).
edge(679, 680).
edge(680, 681).
edge(681, 682).
edge(682, 683).
edge(683, 684).
edge(684, 685).
edge(685, 686).
edge(686, 687).
edge(687, 688).
edge(688, 689).
edge(689, 690).
edge(690, 691).
edge(691, 692).
edge(692, 693).
edge(693, 694).
edge(694, 695).
edge(695, 696).
edge(696, 697).
edge(697, 698).
edge(698, 699).
edge(699, 700).
edge(700, 701).
edge(701, 702).
edge(702, 703).
edge(703, 704).
edge(704, 705).
edge(705, 706).
edge(706, 707).
edge(707, 708).
edge(708, 709).
edge(709, 710).
edge(710, 711).
edge(711, 712).
edge(712, 713).
edge(713, 714).
edge(714, 715).
edge(715, 716).
edge(716, 717).
edge(717, 718).
edge(718, 719).
edge(719, 720).
edge(720, 721).
edge(721, 722).
edge(722, 723).
edge(723, 724).
edge(724, 725).
edge(725, 726).
edge(726, 727).
edge(727, 728).
edge(728, 729).
edge(729, 730).
edge(730, 731).
edge(731, 732).
edge(732, 733).
edge(733, 734).
edge(734, 735).
edge(735, 736).
edge(736, 737).
edge(737, 738).
edge(738, 739).
edge(739, 740).
edge(740, 741).
edge(741, 742).
edge(742, 743).
edge(743, 744).
edge(744, 745).
edge(745, 746).
edge(746, 747).
edge(747, 748).
edge(748, 749).
edge(749, 750).
edge(750, 751).
edge(751, 752).
edge(752, 753).
edge(753, 754).
edge(754, 755).
edge(755, 756).
edge(756, 757).
edge(757, 758).
edge(758, 759).
edge(759, 760).
edge(760, 761).
edge(761, 762).
edge(762, 763).
edge(763, 764).
edge(764, 765).
edge(765, 766).
edge(766, 767).
edge(767, 768).
edge(768, 769).
edge(769, 770).
edge(770, 771).
edge(771, 772).
edge(772, 773).
edge(773, 774).
edge(774, 775).
edge(775, 776).
edge(776, 777).
edge(777, 778).
edge(778, 779).
edge(779, 780).
edge(780, 781).
edge(781, 782).
edge(782, 783).
edge(783, 784).
edge(784, 785).
edge(785, 786).
edge(786, 787).
edge(787, 788).
edge(788, 789).
edge(789, 790).
edge(790, 791).
edge(791, 792).
edge(792, 793).
edge(793, 794).
edge(794, 795).
edge(795, 796).
edge(796, 797).
edge(797, 798).
edge(798, 799).
edge(799, 800).
edge(800, 801).
edge(801, 802).
edge(802, 803).
edge(803, 804).
edge(804, 805).
edge(805, 806).
edge(806, 807).
edge(807, 808).
edge(808, 809).
edge(809, 810).
edge(810, 811).
edge(811, 812).
edge(812, 813).
edge(813, 814).
edge(814, 815).
edge(815, 816).
edge(816, 817).
edge(817, 818).
edge(818, 819).
edge(819, 820).
edge(820, 821).
edge(821, 822).
edge(822, 823).
edge(823, 824).
edge(824, 825).
edge(825, 826).
edge(826, 827).
edge(827, 828).
edge(828, 829).
edge(829, 830).
edge(830, 831).
edge(831, 832).
edge(832, 833).
edge(833, 834).
edge(834, 835).
edge(835, 836).
edge(836, 837).
edge(837, 838).
edge(838, 839).
edge(839, 840).
edge(840, 841).
edge(841, 842).
edge(842, 843).
edge(843, 844).
edge(844, 845).
edge(845, 846).
edge(846, 847).
edge(847, 848).
edge(848, 849).
edge(849, 850).
edge(850, 851).
edge(851, 852).
edge(852, 853).
edge(853, 854).
edge(854, 855).
edge(855, 856).
edge(856, 857).
edge(857, 858).
edge(858, 859).
edge(859, 860).
edge(860, 861).
edge(861, 862).
edge(862, 863).
edge(863, 864).
edge(864, 865).
edge(865, 866).
edge(866, 867).
edge(867, 868).
edge(868, 869).
edge(869, 870).
edge(870, 871).
edge(871, 872).
edge(872, 873).
edge(873, 874).
edge(874, 875).
edge(875, 876).
edge(876, 877).
edge(877, 878).
edge(878, 879).
edge(879, 880).
edge(880, 881).
edge(881, 882).
edge(882, 883).
edge(883, 884).
edge(884, 885).
edge(885, 886).
edge(886, 887).
edge(887, 888).
edge(888, 889).
edge(889, 890).
edge(890, 891).
edge(891, 892).
edge(892, 893).
edge(893, 894).
edge(894, 895).
edge(895, 896).
edge(896, 897).
edge(897, 898).
edge(898, 899).
edge(899, 900).
edge(900, 901).
edge(901, 902).
edge(902, 903).
edge(903, 904).
edge(904, 905).
edge(905, 906).
edge(906, 907).
edge(907, 908).
edge(908, 909).
edge(909, 910).
edge(910, 911).
edge(911, 912).
edge(912, 913).
edge(913, 914).
edge(914, 915).
edge(915, 916).
edge(916, 917).
edge(917, 918).
edge(918, 919).
edge(919, 920).
edge(920, 921).
edge(921, 922).
edge(922, 923).
edge(923, 924).
edge(924, 925).
edge(925, 926).
edge(926, 927).
edge(927, 928).
edge(928, 929).
edge(929, 930).
edge(930, 931).
edge(931, 932).
edge(932, 933).
edge(933, 934).
edge(934, 935).
edge(935, 936).
edge(936, 937).
edge(937, 938).
edge(938, 939).
edge(939, 940).
edge(940, 941).
edge(941, 942).
edge(942, 943).
edge(943, 944).
edge(944, 945).
edge(945, 946).
edge(946, 947).
edge(947, 948).
edge(948, 949).
edge(949, 950).
edge(950, 951).
edge(951, 952).
edge(952, 953).
edge(953, 954).
edge(954, 955).
edge(955, 956).
edge(956, 957).
edge(957, 958).
edge(958, 959).
edge(959, 960).
edge(960, 961).
edge(961, 962).
edge(962, 963).
edge(963, 964).
edge(964, 965).
edge(965, 966).
edge(966, 967).
edge(967, 968).
edge(968, 969).
edge(969, 970).
edge(970, 971).
edge(971, 972).
edge(972, 973).
edge(973, 974).
edge(974, 975).
edge(975, 976).
edge(976, 977).
edge(977, 978).
edge(978, 979).
edge(979, 980).
edge(980, 981).
edge(981, 982).
edge(982, 983).
edge(983, 984).
edge(984, 985).
edge(985, 986).
edge(986, 987).
edge(987, 988).
edge(988, 989).
edge(989, 990).
edge(990, 991).
edge(991, 992).
edge(992, 993).
edge(993, 994).
edge(994, 995).
edge(995, 996).
edge(996, 997).
edge(997, 998).
edge(998, 999).
edge(999, 1000).
edge(1000, 1001).
edge(1001, 1002).
edge(1002, 1003).
edge(1003, 1004).
edge(1004, 1005).
edge(1005, 1006).
edge(1006, 1007).
edge(1007, 1008).
edge(1008, 1009).
edge(1009, 1010).
edge(1010, 1011).
edge(1011, 1012).
edge(1012, 1013).
edge(1013, 1014).
edge(1014, 1015).
edge(1015, 1016).
edge(1016, 1017).
edge(1017, 1018).
edge(1018, 1019).
edge(1019, 1020).
edge(1020, 1021).
edge(1021, 1022).
edge(1022, 1023).
edge(1023, 1024).
edge(1024, 1025).
edge(1025, 1026).
edge(1026, 1027).
edge(1027, 1028).
edge(1028, 1029).
edge(1029, 1030).
edge(1030, 1031).
edge(1031, 1032).
edge(1032, 1033).
edge(1033, 1034).
edge(1034, 1035).
edge(1035, 1036).
edge(1036, 1037).
edge(1037, 1038).
edge(1038, 1039).
edge(1039, 1040).
edge(1040, 1041).
edge(1041, 1042).
edge(1042, 1043).
edge(1043, 1044).
edge(1044, 1045).
edge(1045, 1046).
edge(1046, 1047).
edge(1047, 1048).
edge(1048, 1049).
edge(1049, 1050).
edge(1050, 1051).
edge(1051, 1052).
edge(1052, 1053).
edge(1053, 1054).
edge(1054, 1055).
edge(1055, 1056).
edge(1056, 1057).
edge(1057, 1058).
edge(1058, 1059).
edge(1059, 1060).
edge(1060, 1061).
edge(1061, 1062).
edge(1062, 1063).
edge(1063, 1064).
edge(1064, 1065).
edge(1065, 1066).
edge(1066, 1067).
edge(1067, 1068).
edge(1068, 1069).
edge(1069, 1070).
edge(1070, 1071).
edge(1071, 1072).
edge(1072, 1073).
edge(1073, 1074).
edge(1074, 1075).
edge(1075, 1076).
edge(1076, 1077).
edge(1077, 1078).
edge(1078, 1079).
edge(1079, 1080).
edge(1080, 1081).
edge(1081, 1082).
edge(1082, 1083).
edge(1083, 1084).
edge(1084, 1085).
edge(1085, 1086).
edge(1086, 1087).
edge(1087, 1088).
edge(1088, 1089).
edge(1089, 1090).
edge(1090, 1091).
edge(1091, 1092).
edge(1092, 1093).
edge(1093, 1094).
edge(1094, 1095).
edge(1095, 1096).
edge(1096, 1097).
edge(1097, 1098).
edge(1098, 1099).
edge(1099, 1100).
edge(1100, 1101).
edge(1101, 1102).
edge(1102, 1103).
edge(1103, 1104).
edge(1104, 1105).
edge(1105, 1106).
edge(1106, 1107).
edge(1107, 1108).
edge(1108, 1109).
edge(1109, 1110).
edge(1110, 1111).
edge(1111, 1112).
edge(1112, 1113).
edge(1113, 1114).
edge(1114, 1115).
edge(1115, 1116).
edge(1116, 1117).
edge(1117, 1118).
edge(1118, 1119).
edge(1119, 1120).
edge(1120, 1121).
edge(1121, 1122).
edge(1122, 1123).
edge(1123, 1124).
edge(1124, 1125).
edge(1125, 1126).
edge(1126, 1127).
edge(1127, 1128).
edge(1128, 1129).
edge(1129, 1130).
edge(1130, 1131).
edge(1131, 1132).
edge(1132, 1133).
edge(1133, 1134).
edge(1134, 1135).
edge(1135, 1136).
edge(1136, 1137).
edge(1137, 1138).
edge(1138, 1139).
edge(1139, 1140).
edge(1140, 1141).
edge(1141, 1142).
edge(1142, 1143).
edge(1143, 1144).
edge(1144, 1145).
edge(1145, 1146).
edge(1146, 1147).
edge(1147, 1148).
edge(1148, 1149).
edge(1149, 1150).
edge(1150, 1151).
edge(1151, 1152).
edge(1152, 1153).
edge(1153, 1154).
edge(1154, 1155).
edge(1155, 1156).
edge(1156, 1157).
edge(1157, 1158).
edge(1158, 1159).
edge(1159, 1160).
edge(1160, 1161).
edge(1161, 1162).
edge(1162, 1163).
edge(1163, 1164).
edge(1164, 1165).
edge(1165, 1166).
edge(1166, 1167).
edge(1167, 1168).
edge(1168, 1169).
edge(1169, 1170).
edge(1170, 1171).
edge(1171, 1172).
edge(1172, 1173).
edge(1173, 1174).
edge(1174, 1175).
edge(1175, 1176).
edge(1176, 1177).
edge(1177, 1178).
edge(1178, 1179).
edge(1179, 1180).
edge(1180, 1181).
edge(1181, 1182).
edge(1182, 1183).
edge(1183, 1184).
edge(1184, 1185).
edge(1185, 1186).
edge(1186, 1187).
edge(1187, 1188).
edge(1188, 1189).
edge(1189, 1190).
edge(1190, 1191).
edge(1191, 1192).
edge(1192, 1193).
edge(1193, 1194).
edge(1194, 1195).
edge(1195, 1196).
edge(1196, 1197).
edge(1197, 1198).
edge(1198, 1199).
edge(1199, 1200).
edge(1200, 1201).
edge(1201, 1202).
edge(1202, 1203).
edge(1203, 1204).
edge(1204, 1205).
edge(1205, 1206).
edge(1206, 1207).
edge(1207, 1208).
edge(1208, 1209).
edge(1209, 1210).
edge(1210, 1211).
edge(1211, 1212).
edge(1212, 1213).
edge(1213, 1214).
edge(1214, 1215).
edge(1215, 1216).
edge(1216, 1217).
edge(1217, 1218).
edge(1218, 1219).
edge(1219, 1220).
edge(1220, 1221).
edge(1221, 1222).
edge(1222, 1223).
edge(1223, 1224).
edge(1224, 1225).
edge(1225, 1226).
edge(1226, 1227).
edge(1227, 1228).
edge(1228, 1229).
edge(1229, 1230).
edge(1230, 1231).
edge(1231, 1232).
edge(1232, 1233).
edge(1233, 1234).
edge(1234, 1235).
edge(1235, 1236).
edge(1236, 1237).
edge(1237, 1238).
edge(1238, 1239).
edge(1239, 1240).
edge(1240, 1241).
edge(1241, 1242).
edge(1242, 1243).
edge(1243, 1244).
edge(1244, 1245).
edge(1245, 1246).
edge(1246, 1247).
edge(1247, 1248).
edge(1248, 1249).
edge(1249, 1250).
edge(1250, 1251).
edge(1251, 1252).
edge(1252, 1253).
edge(1253, 1254).
edge(1254, 1255).
edge(1255, 1256).
edge(1256, 1257).
edge(1257, 1258).
edge(1258, 1259).
edge(1259, 1260).
edge(1260, 1261).
edge(1261, 1262).
edge(1262, 1263).
edge(1263, 1264).
edge(1264, 1265).
edge(1265, 1266).
edge(1266, 1267).
edge(1267, 1268).
edge(1268, 1269).
edge(1269, 1270).
edge(1270, 1271).
edge(1271, 1272).
edge(1272, 1273).
edge(1273, 1274).
edge(1274, 1275).
edge(1275, 1276).
edge(1276, 1277).
edge(1277, 1278).
edge(1278, 1279).
edge(1279, 1280).
edge(1280, 1281).
edge(1281, 1282).
edge(1282, 1283).
edge(1283, 1284).
edge(1284, 1285).
edge(1285, 1286).
edge(1286, 1287).
edge(1287, 1288).
edge(1288, 1289).
edge(1289, 1290).
edge(1290, 1291).
edge(1291, 1292).
edge(1292, 1293).
edge(1293, 1294).
edge(1294, 1295).
edge(1295, 1296).
edge(1296, 1297).
edge(1297, 1298).
edge(1298, 1299).
edge(1299, 1300).
edge(1300, 1301).
edge(1301, 1302).
edge(1302, 1303).
edge(1303, 1304).
edge(1304, 1305).
edge(1305, 1306).
edge(1306, 1307).
edge(1307, 1308).
edge(1308, 1309).
edge(1309, 1310).
edge(1310, 1311).
edge(1311, 1312).
edge(1312, 1313).
edge(1313, 1314).
edge(1314, 1315).
edge(1315, 1316).
edge(1316, 1317).
edge(1317, 1318).
edge(1318, 1319).
edge(1319, 1320).
edge(1320, 1321).
edge(1321, 1322).
edge(1322, 1323).
edge(1323, 1324).
edge(1324, 1325).
edge(1325, 1326).
edge(1326, 1327).
edge(1327, 1328).
edge(1328, 1329).
edge(1329, 1330).
edge(1330, 1331).
edge(1331, 1332).
edge(1332, 1333).
edge(1333, 1334).
edge(1334, 1335).
edge(1335, 1336).
edge(1336, 1337).
edge(1337, 1338).
edge(1338, 1339).
edge(1339, 1340).
edge(1340, 1341).
edge(1341, 1342).
edge(1342, 1343).
edge(1343, 1344).
edge(1344, 1345).
edge(1345, 1346).
edge(1346, 1347).
edge(1347, 1348).
edge(1348, 1349).
edge(1349, 1350).
edge(1350, 1351).
edge(1351, 1352).
edge(1352, 1353).
edge(1353, 1354).
edge(1354, 1355).
edge(1355, 1356).
edge(1356, 1357).
edge(1357, 1358).
edge(1358, 1359).
edge(1359, 1360).
edge(1360, 1361).
edge(1361, 1362).
edge(1362, 1363).
edge(1363, 1364).
edge(1364, 1365).
edge(1365, 1366).
edge(1366, 1367).
edge(1367, 1368).
edge(1368, 1369).
edge(1369, 1370).
edge(1370, 1371).
edge(1371, 1372).
edge(1372, 1373).
edge(1373, 1374).
edge(1374, 1375).
edge(1375, 1376).
edge(1376, 1377).
edge(1377, 1378).
edge(1378, 1379).
edge(1379, 1380).
edge(1380, 1381).
edge(1381, 1382).
edge(1382, 1383).
edge(1383, 1384).
edge(1384, 1385).
edge(1385, 1386).
edge(1386, 1387).
edge(1387, 1388).
edge(1388, 1389).
edge(1389, 1390).
edge(1390, 1391).
edge(1391, 1392).
edge(1392, 1393).
edge(1393, 1394).
edge(1394, 1395).
edge(1395, 1396).
edge(1396, 1397).
edge(1397, 1398).
edge(1398, 1399).
edge(1399, 1400).
edge(1400, 1401).
edge(1401, 1402).
edge(1402, 1403).
edge(1403, 1404).
edge(1404, 1405).
edge(1405, 1406).
edge(1406, 1407).
edge(1407, 1408).
edge(1408, 1409).
edge(1409, 1410).
edge(1410, 1411).
edge(1411, 1412).
edge(1412, 1413).
edge(1413, 1414).
edge(1414, 1415).
edge(1415, 1416).
edge(1416, 1417).
edge(1417, 1418).
edge(1418, 1419).
edge(1419, 1420).
edge(1420, 1421).
edge(1421, 1422).
edge(1422, 1423).
edge(1423, 1424).
edge(1424, 1425).
edge(1425, 1426).
edge(1426, 1427).
edge(1427, 1428).
edge(1428, 1429).
edge(1429, 1430).
edge(1430, 1431).
edge(1431, 1432).
edge(1432, 1433).
edge(1433, 1434).
edge(1434, 1435).
edge(1435, 1436).
edge(1436, 1437).
edge(1437, 1438).
edge(1438, 1439).
edge(1439, 1440).
edge(1440, 1441).
edge(1441, 1442).
edge(1442, 1443).
edge(1443, 1444).
edge(1444, 1445).
edge(1445, 1446).
edge(1446, 1447).
edge(1447, 1448).
edge(1448, 1449).
edge(1449, 1450).
edge(1450, 1451).
edge(1451, 1452).
edge(1452, 1453).
edge(1453, 1454).
edge(1454, 1455).
edge(1455, 1456).
edge(1456, 1457).
edge(1457, 1458).
edge(1458, 1459).
edge(1459, 1460).
edge(1460, 1461).
edge(1461, 1462).
edge(1462, 1463).
edge(1463, 1464).
edge(1464, 1465).
edge(1465, 1466).
edge(1466, 1467).
edge(1467, 1468).
edge(1468, 1469).
edge(1469, 1470).
edge(1470, 1471).
edge(1471, 1472).
edge(1472, 1473).
edge(1473, 1474).
edge(1474, 1475).
edge(1475, 1476).
edge(1476, 1477).
edge(1477, 1478).
edge(1478, 1479).
edge(1479, 1480).
edge(1480, 1481).
edge(1481, 1482).
edge(1482, 1483).
edge(1483, 1484).
edge(1484, 1485).
edge(1485, 1486).
edge(1486, 1487).
edge(1487, 1488).
edge(1488, 1489).
edge(1489, 1490).
edge(1490, 1491).
edge(1491, 1492).
edge(1492, 1493).
edge(1493, 1494).
edge(1494, 1495).
edge(1495, 1496).
edge(1496, 1497).
edge(1497, 1498).
edge(1498, 1499).
edge(1499, 1500).
edge(1500, 1501).
edge(1501, 1502).
edge(1502, 1503).
edge(1503, 1504).
edge(1504, 1505).
edge(1505, 1506).
edge(1506, 1507).
edge(1507, 1508).
edge(1508, 1509).
edge(1509, 1510).
edge(1510, 1511).
edge(1511, 1512).
edge(1512, 1513).
edge(1513, 1514).
edge(1514, 1515).
edge(1515, 1516).
edge(1516, 1517).
edge(1517, 1518).
edge(1518, 1519).
edge(1519, 1520).
edge(1520, 1521).
edge(1521, 1522).
edge(1522, 1523).
edge(1523, 1524).
edge(1524, 1525).
edge(1525, 1526).
edge(1526, 1527).
edge(1527, 1528).
edge(1528, 1529).
edge(1529, 1530).
edge(1530, 1531).
edge(1531, 1532).
edge(1532, 1533).
edge(1533, 1534).
edge(1534, 1535).
edge(1535, 1536).
edge(1536, 1537).
edge(1537, 1538).
edge(1538, 1539).
edge(1539, 1540).
edge(1540, 1541).
edge(1541, 1542).
edge(1542, 1543).
edge(1543, 1544).
edge(1544, 1545).
edge(1545, 1546).
edge(1546, 1547).
edge(1547, 1548).
edge(1548, 1549).
edge(1549, 1550).
edge(1550, 1551).
edge(1551, 1552).
edge(1552, 1553).
edge(1553, 1554).
edge(1554, 1555).
edge(1555, 1556).
edge(1556, 1557).
edge(1557, 1558).
edge(1558, 1559).
edge(1559, 1560).
edge(1560, 1561).
edge(1561, 1562).
edge(1562, 1563).
edge(1563, 1564).
edge(1564, 1565).
edge(1565, 1566).
edge(1566, 1567).
edge(1567, 1568).
edge(1568, 1569).
edge(1569, 1570).
edge(1570, 1571).
edge(1571, 1572).
edge(1572, 1573).
edge(1573, 1574).
edge(1574, 1575).
edge(1575, 1576).
edge(1576, 1577).
edge(1577, 1578).
edge(1578, 1579).
edge(1579, 1580).
edge(1580, 1581).
edge(1581, 1582).
edge(1582, 1583).
edge(1583, 1584).
edge(1584, 1585).
edge(1585, 1586).
edge(1586, 1587).
edge(1587, 1588).
edge(1588, 1589).
edge(1589, 1590).
edge(1590, 1591).
edge(1591, 1592).
edge(1592, 1593).
edge(1593, 1594).
edge(1594, 1595).
edge(1595, 1596).
edge(1596, 1597).
edge(1597, 1598).
edge(1598, 1599).
edge(1599, 1600).
edge(1600, 1601).
edge(1601, 1602).
edge(1602, 1603).
edge(1603, 1604).
edge(1604, 1605).
edge(1605, 1606).
edge(1606, 1607).
edge(1607, 1608).
edge(1608, 1609).
edge(1609, 1610).
edge(1610, 1611).
edge(1611, 1612).
edge(1612, 1613).
edge(1613, 1614).
edge(1614, 1615).
edge(1615, 1616).
edge(1616, 1617).
edge(1617, 1618).
edge(1618, 1619).
edge(1619, 1620).
edge(1620, 1621).
edge(1621, 1622).
edge(1622, 1623).
edge(1623, 1624).
edge(1624, 1625).
edge(1625, 1626).
edge(1626, 1627).
edge(1627, 1628).
edge(1628, 1629).
edge(1629, 1630).
edge(1630, 1631).
edge(1631, 1632).
edge(1632, 1633).
edge(1633, 1634).
edge(1634, 1635).
edge(1635, 1636).
edge(1636, 1637).
edge(1637, 1638).
edge(1638, 1639).
edge(1639, 1640).
edge(1640, 1641).
edge(1641, 1642).
edge(1642, 1643).
edge(1643, 1644).
edge(1644, 1645).
edge(1645, 1646).
edge(1646, 1647).
edge(1647, 1648).
edge(1648, 1649).
edge(1649, 1650).
edge(1650, 1651).
edge(1651, 1652).
edge(1652, 1653).
edge(1653, 1654).
edge(1654, 1655).
edge(1655, 1656).
edge(1656, 1657).
edge(1657, 1658).
edge(1658, 1659).
edge(1659, 1660).
edge(1660, 1661).
edge(1661, 1662).
edge(1662, 1663).
edge(1663, 1664).
edge(1664, 1665).
edge(1665, 1666).
edge(1666, 1667).
edge(1667, 1668).
edge(1668, 1669).
edge(1669, 1670).
edge(1670, 1671).
edge(1671, 1672).
edge(1672, 1673).
edge(1673, 1674).
edge(1674, 1675).
edge(1675, 1676).
edge(1676, 1677).
edge(1677, 1678).
edge(1678, 1679).
edge(1679, 1680).
edge(1680, 1681).
edge(1681, 1682).
edge(1682, 1683).
edge(1683, 1684).
edge(1684, 1685).
edge(1685, 1686).
edge(1686, 1687).
edge(1687, 1688).
edge(1688, 1689).
edge(1689, 1690).
edge(1690, 1691).
edge(1691, 1692).
edge(1692, 1693).
edge(1693, 1694).
edge(1694, 1695).
edge(1695, 1696).
edge(1696, 1697).
edge(1697, 1698).
edge(1698, 1699).
edge(1699, 1700).
edge(1700, 1701).
edge(1701, 1702).
edge(1702, 1703).
edge(1703, 1704).
edge(1704, 1705).
edge(1705, 1706).
edge(1706, 1707).
edge(1707, 1708).
edge(1708, 1709).
edge(1709, 1710).
edge(1710, 1711).
edge(1711, 1712).
edge(1712, 1713).
edge(1713, 1714).
edge(1714, 1715).
edge(1715, 1716).
edge(1716, 1717).
edge(1717, 1718).
edge(1718, 1719).
edge(1719, 1720).
edge(1720, 1721).
edge(1721, 1722).
edge(1722, 1723).
edge(1723, 1724).
edge(1724, 1725).
edge(1725, 1726).
edge(1726, 1727).
edge(1727, 1728).
edge(1728, 1729).
edge(1729, 1730).
edge(1730, 1731).
edge(1731, 1732).
edge(1732, 1733).
edge(1733, 1734).
edge(1734, 1735).
edge(1735, 1736).
edge(1736, 1737).
edge(1737, 1738).
edge(1738, 1739).
edge(1739, 1740).
edge(1740, 1741).
edge(1741, 1742).
edge(1742, 1743).
edge(1743, 1744).
edge(1744, 1745).
edge(1745, 1746).
edge(1746, 1747).
edge(1747, 1748).
edge(1748, 1749).
edge(1749, 1750).
edge(1750, 1751).
edge(1751, 1752).
edge(1752, 1753).
edge(1753, 1754).
edge(1754, 1755).
edge(1755, 1756).
edge(1756, 1757).
edge(1757, 1758).
edge(1758, 1759).
edge(1759, 1760).
edge(1760, 1761).
edge(1761, 1762).
edge(1762, 1763).
edge(1763, 1764).
edge(1764, 1765).
edge(1765, 1766).
edge(1766, 1767).
edge(1767, 1768).
edge(1768, 1769).
edge(1769, 1770).
edge(1770, 1771).
edge(1771, 1772).
edge(1772, 1773).
edge(1773, 1774).
edge(1774, 1775).
edge(1775, 1776).
edge(1776, 1777).
edge(1777, 1778).
edge(1778, 1779).
edge(1779, 1780).
edge(1780, 1781).
edge(1781, 1782).
edge(1782, 1783).
edge(1783, 1784).
edge(1784, 1785).
edge(1785, 1786).
edge(1786, 1787).
edge(1787, 1788).
edge(1788, 1789).
edge(1789, 1790).
edge(1790, 1791).
edge(1791, 1792).
edge(1792, 1793).
edge(1793, 1794).
edge(1794, 1795).
edge(1795, 1796).
edge(1796, 1797).
edge(1797, 1798).
edge(1798, 1799).
edge(1799, 1800).
edge(1800, 1801).
edge(1801, 1802).
edge(1802, 1803).
edge(1803, 1804).
edge(1804, 1805).
edge(1805, 1806).
edge(1806, 1807).
edge(1807, 1808).
edge(1808, 1809).
edge(1809, 1810).
edge(1810, 1811).
edge(1811, 1812).
edge(1812, 1813).
edge(1813, 1814).
edge(1814, 1815).
edge(1815, 1816).
edge(1816, 1817).
edge(1817, 1818).
edge(1818, 1819).
edge(1819, 1820).
edge(1820, 1821).
edge(1821, 1822).
edge(1822, 1823).
edge(1823, 1824).
edge(1824, 1825).
edge(1825, 1826).
edge(1826, 1827).
edge(1827, 1828).
edge(1828, 1829).
edge(1829, 1830).
edge(1830, 1831).
edge(1831, 1832).
edge(1832, 1833).
edge(1833, 1834).
edge(1834, 1835).
edge(1835, 1836).
edge(1836, 1837).
edge(1837, 1838).
edge(1838, 1839).
edge(1839, 1840).
edge(1840, 1841).
edge(1841, 1842).
edge(1842, 1843).
edge(1843, 1844).
edge(1844, 1845).
edge(1845, 1846).
edge(1846, 1847).
edge(1847, 1848).
edge(1848, 1849).
edge(1849, 1850).
edge(1850, 1851).
edge(1851, 1852).
edge(1852, 1853).
edge(1853, 1854).
edge(1854, 1855).
edge(1855, 1856).
edge(1856, 1857).
edge(1857, 1858).
edge(1858, 1859).
edge(1859, 1860).
edge(1860, 1861).
edge(1861, 1862).
edge(1862, 1863).
edge(1863, 1864).
edge(1864, 1865).
edge(1865, 1866).
edge(1866, 1867).
edge(1867, 1868).
edge(1868, 1869).
edge(1869, 1870).
edge(1870, 1871).
edge(1871, 1872).
edge(1872, 1873).
edge(1873, 1874).
edge(1874, 1875).
edge(1875, 1876).
edge(1876, 1877).
edge(1877, 1878).
edge(1878, 1879).
edge(1879, 1880).
edge(1880, 1881).
edge(1881, 1882).
edge(1882, 1883).
edge(1883, 1884).
edge(1884, 1885).
edge(1885, 1886).
edge(1886, 1887).
edge(1887, 1888).
edge(1888, 1889).
edge(1889, 1890).
edge(1890, 1891).
edge(1891, 1892).
edge(1892, 1893).
edge(1893, 1894).
edge(1894, 1895).
edge(1895, 1896).
edge(1896, 1897).
edge(1897, 1898).
edge(1898, 1899).
edge(1899, 1900).
edge(1900, 1901).
edge(1901, 1902).
edge(1902, 1903).
edge(1903, 1904).
edge(1904, 1905).
edge(1905, 1906).
edge(1906, 1907).
edge(1907, 1908).
edge(1908, 1909).
edge(1909, 1910).
edge(1910, 1911).
edge(1911, 1912).
edge(1912, 1913).
edge(1913, 1914).
edge(1914, 1915).
edge(1915, 1916).
edge(1916, 1917).
edge(1917, 1918).
edge(1918, 1919).
edge(1919, 1920).
edge(1920, 1921).
edge(1921, 1922).
edge(1922, 1923).
edge(1923, 1924).
edge(1924, 1925).
edge(1925, 1926).
edge(1926, 1927).
edge(1927, 1928).
edge(1928, 1929).
edge(1929, 1930).
edge(1930, 1931).
edge(1931, 1932).
edge(1932, 1933).
edge(1933, 1934).
edge(1934, 1935).
edge(1935, 1936).
edge(1936, 1937).
edge(1937, 1938).
edge(1938, 1939).
edge(1939, 1940).
edge(1940, 1941).
edge(1941, 1942).
edge(1942, 1943).
edge(1943, 1944).
edge(1944, 1945).
edge(1945, 1946).
edge(1946, 1947).
edge(1947, 1948).
edge(1948, 1949).
edge(1949, 1950).
edge(1950, 1951).
edge(1951, 1952).
edge(1952, 1953).
edge(1953, 1954).
edge(1954, 1955).
edge(1955, 1956).
edge(1956, 1957).
edge(1957, 1958).
edge(1958, 1959).
edge(1959, 1960).
edge(1960, 1961).
edge(1961, 1962).
edge(1962, 1963).
edge(1963, 1964).
edge(1964, 1965).
edge(1965, 1966).
edge(1966, 1967).
edge(1967, 1968).
edge(1968, 1969).
edge(1969, 1970).
edge(1970, 1971).
edge(1971, 1972).
edge(1972, 1973).
edge(1973, 1974).
edge(1974, 1975).
edge(1975, 1976).
edge(1976, 1977).
edge(1977, 1978).
edge(1978, 1979).
edge(1979, 1980).
edge(1980, 1981).
edge(1981, 1982).
edge(1982, 1983).
edge(1983, 1984).
edge(1984, 1985).
edge(1985, 1986).
edge(1986, 1987).
edge(1987, 1988).
edge(1988, 1989).
edge(1989, 1990).
edge(1990, 1991).
edge(1991, 1992).
edge(1992, 1993).
edge(1993, 1994).
edge(1994, 1995).
edge(1995, 1996).
edge(1996, 1997).
edge(1997, 1998).
edge(1998, 1999).
edge(1999, 2000).
edge(2000, 2001).
edge(2001, 2002).
edge(2002, 2003).
edge(2003, 2004).
edge(2004, 2005).
edge(2005, 2006).
edge(2006, 2007).
edge(2007, 2008).
edge(2008, 2009).
edge(2009, 2010).
edge(2010, 2011).
edge(2011, 2012).
edge(2012, 2013).
edge(2013, 2014).
edge(2014, 2015).
edge(2015, 2016).
edge(2016, 2017).
edge(2017, 2018).
edge(2018, 2019).
edge(2019, 2020).
edge(2020, 2021).
edge(2021, 2022).
edge(2022, 2023).
edge(2023, 2024).
edge(2024, 2025).
edge(2025, 2026).
edge(2026, 2027).
edge(2027, 2028).
edge(2028, 2029).
edge(2029, 2030).
edge(2030, 2031).
edge(2031, 2032).
edge(2032, 2033).
edge(2033, 2034).
edge(2034, 2035).
edge(2035, 2036).
edge(2036, 2037).
edge(2037, 2038).
edge(2038, 2039).
edge(2039, 2040).
edge(2040, 2041).
edge(2041, 2042).
edge(2042, 2043).
edge(2043, 2044).
edge(2044, 2045).
edge(2045, 2046).
edge(2046, 2047).
edge(2047, 2048).
edge(2048, 2049).
edge(2049, 2050).
edge(2050, 2051).
edge(2051, 2052).
edge(2052, 2053).
edge(2053, 2054).
edge(2054, 2055).
edge(2055, 2056).
edge(2056, 2057).
edge(2057, 2058).
edge(2058, 2059).
edge(2059, 2060).
edge(2060, 2061).
edge(2061, 2062).
edge(2062, 2063).
edge(2063, 2064).
edge(2064, 2065).
edge(2065, 2066).
edge(2066, 2067).
edge(2067, 2068).
edge(2068, 2069).
edge(2069, 2070).
edge(2070, 2071).
edge(2071, 2072).
edge(2072, 2073).
edge(2073, 2074).
edge(2074, 2075).
edge(2075, 2076).
edge(2076, 2077).
edge(2077, 2078).
edge(2078, 2079).
edge(2079, 2080).
edge(2080, 2081).
edge(2081, 2082).
edge(2082, 2083).
edge(2083, 2084).
edge(2084, 2085).
edge(2085, 2086).
edge(2086, 2087).
edge(2087, 2088).
edge(2088, 2089).
edge(2089, 2090).
edge(2090, 2091).
edge(2091, 2092).
edge(2092, 2093).
edge(2093, 2094).
edge(2094, 2095).
edge(2095, 2096).
edge(2096, 2097).
edge(2097, 2098).
edge(2098, 2099).
edge(2099, 2100).
edge(2100, 2101).
edge(2101, 2102).
edge(2102, 2103).
edge(2103, 2104).
edge(2104, 2105).
edge(2105, 2106).
edge(2106, 2107).
edge(2107, 2108).
edge(2108, 2109).
edge(2109, 2110).
edge(2110, 2111).
edge(2111, 2112).
edge(2112, 2113).
edge(2113, 2114).
edge(2114, 2115).
edge(2115, 2116).
edge(2116, 2117).
edge(2117, 2118).
edge(2118, 2119).
edge(2119, 2120).
edge(2120, 2121).
edge(2121, 2122).
edge(2122, 2123).
edge(2123, 2124).
edge(2124, 2125).
edge(2125, 2126).
edge(2126, 2127).
edge(2127, 2128).
edge(2128, 2129).
edge(2129, 2130).
edge(2130, 2131).
edge(2131, 2132).
edge(2132, 2133).
edge(2133, 2134).
edge(2134, 2135).
edge(2135, 2136).
edge(2136, 2137).
edge(2137, 2138).
edge(2138, 2139).
edge(2139, 2140).
edge(2140, 2141).
edge(2141, 2142).
edge(2142, 2143).
edge(2143, 2144).
edge(2144, 2145).
edge(2145, 2146).
edge(2146, 2147).
edge(2147, 2148).
edge(2148, 2149).
edge(2149, 2150).
edge(2150, 2151).
edge(2151, 2152).
edge(2152, 2153).
edge(2153, 2154).
edge(2154, 2155).
edge(2155, 2156).
edge(2156, 2157).
edge(2157, 2158).
edge(2158, 2159).
edge(2159, 2160).
edge(2160, 2161).
edge(2161, 2162).
edge(2162, 2163).
edge(2163, 2164).
edge(2164, 2165).
edge(2165, 2166).
edge(2166, 2167).
edge(2167, 2168).
edge(2168, 2169).
edge(2169, 2170).
edge(2170, 2171).
edge(2171, 2172).
edge(2172, 2173).
edge(2173, 2174).
edge(2174, 2175).
edge(2175, 2176).
edge(2176, 2177).
edge(2177, 2178).
edge(2178, 2179).
edge(2179, 2180).
edge(2180, 2181).
edge(2181, 2182).
edge(2182, 2183).
edge(2183, 2184).
edge(2184, 2185).
edge(2185, 2186).
edge(2186, 2187).
edge(2187, 2188).
edge(2188, 2189).
edge(2189, 2190).
edge(2190, 2191).
edge(2191, 2192).
edge(2192, 2193).
edge(2193, 2194).
edge(2194, 2195).
edge(2195, 2196).
edge(2196, 2197).
edge(2197, 2198).
edge(2198, 2199).
edge(2199, 2200).
edge(2200, 2201).
edge(2201, 2202).
edge(2202, 2203).
edge(2203, 2204).
edge(2204, 2205).
edge(2205, 2206).
edge(2206, 2207).
edge(2207, 2208).
edge(2208, 2209).
edge(2209, 2210).
edge(2210, 2211).
edge(2211, 2212).
edge(2212, 2213).
edge(2213, 2214).
edge(2214, 2215).
edge(2215, 2216).
edge(2216, 2217).
edge(2217, 2218).
edge(2218, 2219).
edge(2219, 2220).
edge(2220, 2221).
edge(2221, 2222).
edge(2222, 2223).
edge(2223, 2224).
edge(2224, 2225).
edge(2225, 2226).
edge(2226, 2227).
edge(2227, 2228).
edge(2228, 2229).
edge(2229, 2230).
edge(2230, 2231).
edge(2231, 2232).
edge(2232, 2233).
edge(2233, 2234).
edge(2234, 2235).
edge(2235, 2236).
edge(2236, 2237).
edge(2237, 2238).
edge(2238, 2239).
edge(2239, 2240).
edge(2240, 2241).
edge(2241, 2242).
edge(2242, 2243).
edge(2243, 2244).
edge(2244, 2245).
edge(2245, 2246).
edge(2246, 2247).
edge(2247, 2248).
edge(2248, 2249).
edge(2249, 2250).
edge(2250, 2251).
edge(2251, 2252).
edge(2252, 2253).
edge(2253, 2254).
edge(2254, 2255).
edge(2255, 2256).
edge(2256, 2257).
edge(2257, 2258).
edge(2258, 2259).
edge(2259, 2260).
edge(2260, 2261).
edge(2261, 2262).
edge(2262, 2263).
edge(2263, 2264).
edge(2264, 2265).
edge(2265, 2266).
edge(2266, 2267).
edge(2267, 2268).
edge(2268, 2269).
edge(2269, 2270).
edge(2270, 2271).
edge(2271, 2272).
edge(2272, 2273).
edge(2273, 2274).
edge(2274, 2275).
edge(2275, 2276).
edge(2276, 2277).
edge(2277, 2278).
edge(2278, 2279).
edge(2279, 2280).
edge(2280, 2281).
edge(2281, 2282).
edge(2282, 2283).
edge(2283, 2284).
edge(2284, 2285).
edge(2285, 2286).
edge(2286, 2287).
edge(2287, 2288).
edge(2288, 2289).
edge(2289, 2290).
edge(2290, 2291).
edge(2291, 2292).
edge(2292, 2293).
edge(2293, 2294).
edge(2294, 2295).
edge(2295, 2296).
edge(2296, 2297).
edge(2297, 2298).
edge(2298, 2299).
edge(2299, 2300).
edge(2300, 2301).
edge(2301, 2302).
edge(2302, 2303).
edge(2303, 2304).
edge(2304, 2305).
edge(2305, 2306).
edge(2306, 2307).
edge(2307, 2308).
edge(2308, 2309).
edge(2309, 2310).
edge(2310, 2311).
edge(2311, 2312).
edge(2312, 2313).
edge(2313, 2314).
edge(2314, 2315).
edge(2315, 2316).
edge(2316, 2317).
edge(2317, 2318).
edge(2318, 2319).
edge(2319, 2320).
edge(2320, 2321).
edge(2321, 2322).
edge(2322, 2323).
edge(2323, 2324).
edge(2324, 2325).
edge(2325, 2326).
edge(2326, 2327).
edge(2327, 2328).
edge(2328, 2329).
edge(2329, 2330).
edge(2330, 2331).
edge(2331, 2332).
edge(2332, 2333).
edge(2333, 2334).
edge(2334, 2335).
edge(2335, 2336).
edge(2336, 2337).
edge(2337, 2338).
edge(2338, 2339).
edge(2339, 2340).
edge(2340, 2341).
edge(2341, 2342).
edge(2342, 2343).
edge(2343, 2344).
edge(2344, 2345).
edge(2345, 2346).
edge(2346, 2347).
edge(2347, 2348).
edge(2348, 2349).
edge(2349, 2350).
edge(2350, 2351).
edge(2351, 2352).
edge(2352, 2353).
edge(2353, 2354).
edge(2354, 2355).
edge(2355, 2356).
edge(2356, 2357).
edge(2357, 2358).
edge(2358, 2359).
edge(2359, 2360).
edge(2360, 2361).
edge(2361, 2362).
edge(2362, 2363).
edge(2363, 2364).
edge(2364, 2365).
edge(2365, 2366).
edge(2366, 2367).
edge(2367, 2368).
edge(2368, 2369).
edge(2369, 2370).
edge(2370, 2371).
edge(2371, 2372).
edge(2372, 2373).
edge(2373, 2374).
edge(2374, 2375).
edge(2375, 2376).
edge(2376, 2377).
edge(2377, 2378).
edge(2378, 2379).
edge(2379, 2380).
edge(2380, 2381).
edge(2381, 2382).
edge(2382, 2383).
edge(2383, 2384).
edge(2384, 2385).
edge(2385, 2386).
edge(2386, 2387).
edge(2387, 2388).
edge(2388, 2389).
edge(2389, 2390).
edge(2390, 2391).
edge(2391, 2392).
edge(2392, 2393).
edge(2393, 2394).
edge(2394, 2395).
edge(2395, 2396).
edge(2396, 2397).
edge(2397, 2398).
edge(2398, 2399).
edge(2399, 2400).
edge(2400, 2401).
edge(2401, 2402).
edge(2402, 2403).
edge(2403, 2404).
edge(2404, 2405).
edge(2405, 2406).
edge(2406, 2407).
edge(2407, 2408).
edge(2408, 2409).
edge(2409, 2410).
edge(2410, 2411).
edge(2411, 2412).
edge(2412, 2413).
edge(2413, 2414).
edge(2414, 2415).
edge(2415, 2416).
edge(2416, 2417).
edge(2417, 2418).
edge(2418, 2419).
edge(2419, 2420).
edge(2420, 2421).
edge(2421, 2422).
edge(2422, 2423).
edge(2423, 2424).
edge(2424, 2425).
edge(2425, 2426).
edge(2426, 2427).
edge(2427, 2428).
edge(2428, 2429).
edge(2429, 2430).
edge(2430, 2431).
edge(2431, 2432).
edge(2432, 2433).
edge(2433, 2434).
edge(2434, 2435).
edge(2435, 2436).
edge(2436, 2437).
edge(2437, 2438).
edge(2438, 2439).
edge(2439, 2440).
edge(2440, 2441).
edge(2441, 2442).
edge(2442, 2443).
edge(2443, 2444).
edge(2444, 2445).
edge(2445, 2446).
edge(2446, 2447).
edge(2447, 2448).
edge(2448, 2449).
edge(2449, 2450).
edge(2450, 2451).
edge(2451, 2452).
edge(2452, 2453).
edge(2453, 2454).
edge(2454, 2455).
edge(2455, 2456).
edge(2456, 2457).
edge(2457, 2458).
edge(2458, 2459).
edge(2459, 2460).
edge(2460, 2461).
edge(2461, 2462).
edge(2462, 2463).
edge(2463, 2464).
edge(2464, 2465).
edge(2465, 2466).
edge(2466, 2467).
edge(2467, 2468).
edge(2468, 2469).
edge(2469, 2470).
edge(2470, 2471).
edge(2471, 2472).
edge(2472, 2473).
edge(2473, 2474).
edge(2474, 2475).
edge(2475, 2476).
edge(2476, 2477).
edge(2477, 2478).
edge(2478, 2479).
edge(2479, 2480).
edge(2480, 2481).
edge(2481, 2482).
edge(2482, 2483).
edge(2483, 2484).
edge(2484, 2485).
edge(2485, 2486).
edge(2486, 2487).
edge(2487, 2488).
edge(2488, 2489).
edge(2489, 2490).
edge(2490, 2491).
edge(2491, 2492).
edge(2492, 2493).
edge(2493, 2494).
edge(2494, 2495).
edge(2495, 2496).
edge(2496, 2497).
edge(2497, 2498).
edge(2498, 2499).
edge(2499, 2500).
edge(2500, 2501).
edge(2501, 2502).
edge(2502, 2503).
edge(2503, 2504).
edge(2504, 2505).
edge(2505, 2506).
edge(2506, 2507).
edge(2507, 2508).
edge(2508, 2509).
edge(2509, 2510).
edge(2510, 2511).
edge(2511, 2512).
edge(2512, 2513).
edge(2513, 2514).
edge(2514, 2515).
edge(2515, 2516).
edge(2516, 2517).
edge(2517, 2518).
edge(2518, 2519).
edge(2519, 2520).
edge(2520, 2521).
edge(2521, 2522).
edge(2522, 2523).
edge(2523, 2524).
edge(2524, 2525).
edge(2525, 2526).
edge(2526, 2527).
edge(2527, 2528).
edge(2528, 2529).
edge(2529, 2530).
edge(2530, 2531).
edge(2531, 2532).
edge(2532, 2533).
edge(2533, 2534).
edge(2534, 2535).
edge(2535, 2536).
edge(2536, 2537).
edge(2537, 2538).
edge(2538, 2539).
edge(2539, 2540).
edge(2540, 2541).
edge(2541, 2542).
edge(2542, 2543).
edge(2543, 2544).
edge(2544, 2545).
edge(2545, 2546).
edge(2546, 2547).
edge(2547, 2548).
edge(2548, 2549).
edge(2549, 2550).
edge(2550, 2551).
edge(2551, 2552).
edge(2552, 2553).
edge(2553, 2554).
edge(2554, 2555).
edge(2555, 2556).
edge(2556, 2557).
edge(2557, 2558).
edge(2558, 2559).
edge(2559, 2560).
edge(2560, 2561).
edge(2561, 2562).
edge(2562, 2563).
edge(2563, 2564).
edge(2564, 2565).
edge(2565, 2566).
edge(2566, 2567).
edge(2567, 2568).
edge(2568, 2569).
edge(2569, 2570).
edge(2570, 2571).
edge(2571, 2572).
edge(2572, 2573).
edge(2573, 2574).
edge(2574, 2575).
edge(2575, 2576).
edge(2576, 2577).
edge(2577, 2578).
edge(2578, 2579).
edge(2579, 2580).
edge(2580, 2581).
edge(2581, 2582).
edge(2582, 2583).
edge(2583, 2584).
edge(2584, 2585).
edge(2585, 2586).
edge(2586, 2587).
edge(2587, 2588).
edge(2588, 2589).
edge(2589, 2590).
edge(2590, 2591).
edge(2591, 2592).
edge(2592, 2593).
edge(2593, 2594).
edge(2594, 2595).
edge(2595, 2596).
edge(2596, 2597).
edge(2597, 2598).
edge(2598, 2599).
edge(2599, 2600).
edge(2600, 2601).
edge(2601, 2602).
edge(2602, 2603).
edge(2603, 2604).
edge(2604, 2605).
edge(2605, 2606).
edge(2606, 2607).
edge(2607, 2608).
edge(2608, 2609).
edge(2609, 2610).
edge(2610, 2611).
edge(2611, 2612).
edge(2612, 2613).
edge(2613, 2614).
edge(2614, 2615).
edge(2615, 2616).
edge(2616, 2617).
edge(2617, 2618).
edge(2618, 2619).
edge(2619, 2620).
edge(2620, 2621).
edge(2621, 2622).
edge(2622, 2623).
edge(2623, 2624).
edge(2624, 2625).
edge(2625, 2626).
edge(2626, 2627).
edge(2627, 2628).
edge(2628, 2629).
edge(2629, 2630).
edge(2630, 2631).
edge(2631, 2632).
edge(2632, 2633).
edge(2633, 2634).
edge(2634, 2635).
edge(2635, 2636).
edge(2636, 2637).
edge(2637, 2638).
edge(2638, 2639).
edge(2639, 2640).
edge(2640, 2641).
edge(2641, 2642).
edge(2642, 2643).
edge(2643, 2644).
edge(2644, 2645).
edge(2645, 2646).
edge(2646, 2647).
edge(2647, 2648).
edge(2648, 2649).
edge(2649, 2650).
edge(2650, 2651).
edge(2651, 2652).
edge(2652, 2653).
edge(2653, 2654).
edge(2654, 2655).
edge(2655, 2656).
edge(2656, 2657).
edge(2657, 2658).
edge(2658, 2659).
edge(2659, 2660).
edge(2660, 2661).
edge(2661, 2662).
edge(2662, 2663).
edge(2663, 2664).
edge(2664, 2665).
edge(2665, 2666).
edge(2666, 2667).
edge(2667, 2668).
edge(2668, 2669).
edge(2669, 2670).
edge(2670, 2671).
edge(2671, 2672).
edge(2672, 2673).
edge(2673, 2674).
edge(2674, 2675).
edge(2675, 2676).
edge(2676, 2677).
edge(2677, 2678).
edge(2678, 2679).
edge(2679, 2680).
edge(2680, 2681).
edge(2681, 2682).
edge(2682, 2683).
edge(2683, 2684).
edge(2684, 2685).
edge(2685, 2686).
edge(2686, 2687).
edge(2687, 2688).
edge(2688, 2689).
edge(2689, 2690).
edge(2690, 2691).
edge(2691, 2692).
edge(2692, 2693).
edge(2693, 2694).
edge(2694, 2695).
edge(2695, 2696).
edge(2696, 2697).
edge(2697, 2698).
edge(2698, 2699).
edge(2699, 2700).
edge(2700, 2701).
edge(2701, 2702).
edge(2702, 2703).
edge(2703, 2704).
edge(2704, 2705).
edge(2705, 2706).
edge(2706, 2707).
edge(2707, 2708).
edge(2708, 2709).
edge(2709, 2710).
edge(2710, 2711).
edge(2711, 2712).
edge(2712, 2713).
edge(2713, 2714).
edge(2714, 2715).
edge(2715, 2716).
edge(2716, 2717).
edge(2717, 2718).
edge(2718, 2719).
edge(2719, 2720).
edge(2720, 2721).
edge(2721, 2722).
edge(2722, 2723).
edge(2723, 2724).
edge(2724, 2725).
edge(2725, 2726).
edge(2726, 2727).
edge(2727, 2728).
edge(2728, 2729).
edge(2729, 2730).
edge(2730, 2731).
edge(2731, 2732).
edge(2732, 2733).
edge(2733, 2734).
edge(2734, 2735).
edge(2735, 2736).
edge(2736, 2737).
edge(2737, 2738).
edge(2738, 2739).
edge(2739, 2740).
edge(2740, 2741).
edge(2741, 2742).
edge(2742, 2743).
edge(2743, 2744).
edge(2744, 2745).
edge(2745, 2746).
edge(2746, 2747).
edge(2747, 2748).
edge(2748, 2749).
edge(2749, 2750).
edge(2750, 2751).
edge(2751, 2752).
edge(2752, 2753).
edge(2753, 2754).
edge(2754, 2755).
edge(2755, 2756).
edge(2756, 2757).
edge(2757, 2758).
edge(2758, 2759).
edge(2759, 2760).
edge(2760, 2761).
edge(2761, 2762).
edge(2762, 2763).
edge(2763, 2764).
edge(2764, 2765).
edge(2765, 2766).
edge(2766, 2767).
edge(2767, 2768).
edge(2768, 2769).
edge(2769, 2770).
edge(2770, 2771).
edge(2771, 2772).
edge(2772, 2773).
edge(2773, 2774).
edge(2774, 2775).
edge(2775, 2776).
edge(2776, 2777).
edge(2777, 2778).
edge(2778, 2779).
edge(2779, 2780).
edge(2780, 2781).
edge(2781, 2782).
edge(2782, 2783).
edge(2783, 2784).
edge(2784, 2785).
edge(2785, 2786).
edge(2786, 2787).
edge(2787, 2788).
edge(2788, 2789).
edge(2789, 2790).
edge(2790, 2791).
edge(2791, 2792).
edge(2792, 2793).
edge(2793, 2794).
edge(2794, 2795).
edge(2795, 2796).
edge(2796, 2797).
edge(2797, 2798).
edge(2798, 2799).
edge(2799, 2800).
edge(2800, 2801).
edge(2801, 2802).
edge(2802, 2803).
edge(2803, 2804).
edge(2804, 2805).
edge(2805, 2806).
edge(2806, 2807).
edge(2807, 2808).
edge(2808, 2809).
edge(2809, 2810).
edge(2810, 2811).
edge(2811, 2812).
edge(2812, 2813).
edge(2813, 2814).
edge(2814, 2815).
edge(2815, 2816).
edge(2816, 2817).
edge(2817, 2818).
edge(2818, 2819).
edge(2819, 2820).
edge(2820, 2821).
edge(2821, 2822).
edge(2822, 2823).
edge(2823, 2824).
edge(2824, 2825).
edge(2825, 2826).
edge(2826, 2827).
edge(2827, 2828).
edge(2828, 2829).
edge(2829, 2830).
edge(2830, 2831).
edge(2831, 2832).
edge(2832, 2833).
edge(2833, 2834).
edge(2834, 2835).
edge(2835, 2836).
edge(2836, 2837).
edge(2837, 2838).
edge(2838, 2839).
edge(2839, 2840).
edge(2840, 2841).
edge(2841, 2842).
edge(2842, 2843).
edge(2843, 2844).
edge(2844, 2845).
edge(2845, 2846).
edge(2846, 2847).
edge(2847, 2848).
edge(2848, 2849).
edge(2849, 2850).
edge(2850, 2851).
edge(2851, 2852).
edge(2852, 2853).
edge(2853, 2854).
edge(2854, 2855).
edge(2855, 2856).
edge(2856, 2857).
edge(2857, 2858).
edge(2858, 2859).
edge(2859, 2860).
edge(2860, 2861).
edge(2861, 2862).
edge(2862, 2863).
edge(2863, 2864).
edge(2864, 2865).
edge(2865, 2866).
edge(2866, 2867).
edge(2867, 2868).
edge(2868, 2869).
edge(2869, 2870).
edge(2870, 2871).
edge(2871, 2872).
edge(2872, 2873).
edge(2873, 2874).
edge(2874, 2875).
edge(2875, 2876).
edge(2876, 2877).
edge(2877, 2878).
edge(2878, 2879).
edge(2879, 2880).
edge(2880, 2881).
edge(2881, 2882).
edge(2882, 2883).
edge(2883, 2884).
edge(2884, 2885).
edge(2885, 2886).
edge(2886, 2887).
edge(2887, 2888).
edge(2888, 2889).
edge(2889, 2890).
edge(2890, 2891).
edge(2891, 2892).
edge(2892, 2893).
edge(2893, 2894).
edge(2894, 2895).
edge(2895, 2896).
edge(2896, 2897).
edge(2897, 2898).
edge(2898, 2899).
edge(2899, 2900).
edge(2900, 2901).
edge(2901, 2902).
edge(2902, 2903).
edge(2903, 2904).
edge(2904, 2905).
edge(2905, 2906).
edge(2906, 2907).
edge(2907, 2908).
edge(2908, 2909).
edge(2909, 2910).
edge(2910, 2911).
edge(2911, 2912).
edge(2912, 2913).
edge(2913, 2914).
edge(2914, 2915).
edge(2915, 2916).
edge(2916, 2917).
edge(2917, 2918).
edge(2918, 2919).
edge(2919, 2920).
edge(2920, 2921).
edge(2921, 2922).
edge(2922, 2923).
edge(2923, 2924).
edge(2924, 2925).
edge(2925, 2926).
edge(2926, 2927).
edge(2927, 2928).
edge(2928, 2929).
edge(2929, 2930).
edge(2930, 2931).
edge(2931, 2932).
edge(2932, 2933).
edge(2933, 2934).
edge(2934, 2935).
edge(2935, 2936).
edge(2936, 2937).
edge(2937, 2938).
edge(2938, 2939).
edge(2939, 2940).
edge(2940, 2941).
edge(2941, 2942).
edge(2942, 2943).
edge(2943, 2944).
edge(2944, 2945).
edge(2945, 2946).
edge(2946, 2947).
edge(2947, 2948).
edge(2948, 2949).
edge(2949, 2950).
edge(2950, 2951).
edge(2951, 2952).
edge(2952, 2953).
edge(2953, 2954).
edge(2954, 2955).
edge(2955, 2956).
edge(2956, 2957).
edge(2957, 2958).
edge(2958, 2959).
edge(2959, 2960).
edge(2960, 2961).
edge(2961, 2962).
edge(2962, 2963).
edge(2963, 2964).
edge(2964, 2965).
edge(2965, 2966).
edge(2966, 2967).
edge(2967, 2968).
edge(2968, 2969).
edge(2969, 2970).
edge(2970, 2971).
edge(2971, 2972).
edge(2972, 2973).
edge(2973, 2974).
edge(2974, 2975).
edge(2975, 2976).
edge(2976, 2977).
edge(2977, 2978).
edge(2978, 2979).
edge(2979, 2980).
edge(2980, 2981).
edge(2981, 2982).
edge(2982, 2983).
edge(2983, 2984).
edge(2984, 2985).
edge(2985, 2986).
edge(2986, 2987).
edge(2987, 2988).
edge(2988, 2989).
edge(2989, 2990).
edge(2990, 2991).
edge(2991, 2992).
edge(2992, 2993).
edge(2993, 2994).
edge(2994, 2995).
edge(2995, 2996).
edge(2996, 2997).
edge(2997, 2998).
edge(2998, 2999).
edge(2999, 3000).
edge(3000, 3001).
edge(3001, 3002).
edge(3002, 3003).
edge(3003, 3004).
edge(3004, 3005).
edge(3005, 3006).
edge(3006, 3007).
edge(3007, 3008).
edge(3008, 3009).
edge(3009, 3010).
edge(3010, 3011).
edge(3011, 3012).
edge(3012, 3013).
edge(3013, 3014).
edge(3014, 3015).
edge(3015, 3016).
edge(3016, 3017).
edge(3017, 3018).
edge(3018, 3019).
edge(3019, 3020).
edge(3020, 3021).
edge(3021, 3022).
edge(3022, 3023).
edge(3023, 3024).
edge(3024, 3025).
edge(3025, 3026).
edge(3026, 3027).
edge(3027, 3028).
edge(3028, 3029).
edge(3029, 3030).
edge(3030, 3031).
edge(3031, 3032).
edge(3032, 3033).
edge(3033, 3034).
edge(3034, 3035).
edge(3035, 3036).
edge(3036, 3037).
edge(3037, 3038).
edge(3038, 3039).
edge(3039, 3040).
edge(3040, 3041).
edge(3041, 3042).
edge(3042, 3043).
edge(3043, 3044).
edge(3044, 3045).
edge(3045, 3046).
edge(3046, 3047).
edge(3047, 3048).
edge(3048, 3049).
edge(3049, 3050).
edge(3050, 3051).
edge(3051, 3052).
edge(3052, 3053).
edge(3053, 3054).
edge(3054, 3055).
edge(3055, 3056).
edge(3056, 3057).
edge(3057, 3058).
edge(3058, 3059).
edge(3059, 3060).
edge(3060, 3061).
edge(3061, 3062).
edge(3062, 3063).
edge(3063, 3064).
edge(3064, 3065).
edge(3065, 3066).
edge(3066, 3067).
edge(3067, 3068).
edge(3068, 3069).
edge(3069, 3070).
edge(3070, 3071).
edge(3071, 3072).
edge(3072, 3073).
edge(3073, 3074).
edge(3074, 3075).
edge(3075, 3076).
edge(3076, 3077).
edge(3077, 3078).
edge(3078, 3079).
edge(3079, 3080).
edge(3080, 3081).
edge(3081, 3082).
edge(3082, 3083).
edge(3083, 3084).
edge(3084, 3085).
edge(3085, 3086).
edge(3086, 3087).
edge(3087, 3088).
edge(3088, 3089).
edge(3089, 3090).
edge(3090, 3091).
edge(3091, 3092).
edge(3092, 3093).
edge(3093, 3094).
edge(3094, 3095).
edge(3095, 3096).
edge(3096, 3097).
edge(3097, 3098).
edge(3098, 3099).
edge(3099, 3100).
edge(3100, 3101).
edge(3101, 3102).
edge(3102, 3103).
edge(3103, 3104).
edge(3104, 3105).
edge(3105, 3106).
edge(3106, 3107).
edge(3107, 3108).
edge(3108, 3109).
edge(3109, 3110).
edge(3110, 3111).
edge(3111, 3112).
edge(3112, 3113).
edge(3113, 3114).
edge(3114, 3115).
edge(3115, 3116).
edge(3116, 3117).
edge(3117, 3118).
edge(3118, 3119).
edge(3119, 3120).
edge(3120, 3121).
edge(3121, 3122).
edge(3122, 3123).
edge(3123, 3124).
edge(3124, 3125).
edge(3125, 3126).
edge(3126, 3127).
edge(3127, 3128).
edge(3128, 3129).
edge(3129, 3130).
edge(3130, 3131).
edge(3131, 3132).
edge(3132, 3133).
edge(3133, 3134).
edge(3134, 3135).
edge(3135, 3136).
edge(3136, 3137).
edge(3137, 3138).
edge(3138, 3139).
edge(3139, 3140).
edge(3140, 3141).
edge(3141, 3142).
edge(3142, 3143).
edge(3143, 3144).
edge(3144, 3145).
edge(3145, 3146).
edge(3146, 3147).
edge(3147, 3148).
edge(3148, 3149).
edge(3149, 3150).
edge(3150, 3151).
edge(3151, 3152).
edge(3152, 3153).
edge(3153, 3154).
edge(3154, 3155).
edge(3155, 3156).
edge(3156, 3157).
edge(3157, 3158).
edge(3158, 3159).
edge(3159, 3160).
edge(3160, 3161).
edge(3161, 3162).
edge(3162, 3163).
edge(3163, 3164).
edge(3164, 3165).
edge(3165, 3166).
edge(3166, 3167).
edge(3167, 3168).
edge(3168, 3169).
edge(3169, 3170).
edge(3170, 3171).
edge(3171, 3172).
edge(3172, 3173).
edge(3173, 3174).
edge(3174, 3175).
edge(3175, 3176).
edge(3176, 3177).
edge(3177, 3178).
edge(3178, 3179).
edge(3179, 3180).
edge(3180, 3181).
edge(3181, 3182).
edge(3182, 3183).
edge(3183, 3184).
edge(3184, 3185).
edge(3185, 3186).
edge(3186, 3187).
edge(3187, 3188).
edge(3188, 3189).
edge(3189, 3190).
edge(3190, 3191).
edge(3191, 3192).
edge(3192, 3193).
edge(3193, 3194).
edge(3194, 3195).
edge(3195, 3196).
edge(3196, 3197).
edge(3197, 3198).
edge(3198, 3199).
edge(3199, 3200).
edge(3200, 3201).
edge(3201, 3202).
edge(3202, 3203).
edge(3203, 3204).
edge(3204, 3205).
edge(3205, 3206).
edge(3206, 3207).
edge(3207, 3208).
edge(3208, 3209).
edge(3209, 3210).
edge(3210, 3211).
edge(3211, 3212).
edge(3212, 3213).
edge(3213, 3214).
edge(3214, 3215).
edge(3215, 3216).
edge(3216, 3217).
edge(3217, 3218).
edge(3218, 3219).
edge(3219, 3220).
edge(3220, 3221).
edge(3221, 3222).
edge(3222, 3223).
edge(3223, 3224).
edge(3224, 3225).
edge(3225, 3226).
edge(3226, 3227).
edge(3227, 3228).
edge(3228, 3229).
edge(3229, 3230).
edge(3230, 3231).
edge(3231, 3232).
edge(3232, 3233).
edge(3233, 3234).
edge(3234, 3235).
edge(3235, 3236).
edge(3236, 3237).
edge(3237, 3238).
edge(3238, 3239).
edge(3239, 3240).
edge(3240, 3241).
edge(3241, 3242).
edge(3242, 3243).
edge(3243, 3244).
edge(3244, 3245).
edge(3245, 3246).
edge(3246, 3247).
edge(3247, 3248).
edge(3248, 3249).
edge(3249, 3250).
edge(3250, 3251).
edge(3251, 3252).
edge(3252, 3253).
edge(3253, 3254).
edge(3254, 3255).
edge(3255, 3256).
edge(3256, 3257).
edge(3257, 3258).
edge(3258, 3259).
edge(3259, 3260).
edge(3260, 3261).
edge(3261, 3262).
edge(3262, 3263).
edge(3263, 3264).
edge(3264, 3265).
edge(3265, 3266).
edge(3266, 3267).
edge(3267, 3268).
edge(3268, 3269).
edge(3269, 3270).
edge(3270, 3271).
edge(3271, 3272).
edge(3272, 3273).
edge(3273, 3274).
edge(3274, 3275).
edge(3275, 3276).
edge(3276, 3277).
edge(3277, 3278).
edge(3278, 3279).
edge(3279, 3280).
edge(3280, 3281).
edge(3281, 3282).
edge(3282, 3283).
edge(3283, 3284).
edge(3284, 3285).
edge(3285, 3286).
edge(3286, 3287).
edge(3287, 3288).
edge(3288, 3289).
edge(3289, 3290).
edge(3290, 3291).
edge(3291, 3292).
edge(3292, 3293).
edge(3293, 3294).
edge(3294, 3295).
edge(3295, 3296).
edge(3296, 3297).
edge(3297, 3298).
edge(3298, 3299).
edge(3299, 3300).
edge(3300, 3301).
edge(3301, 3302).
edge(3302, 3303).
edge(3303, 3304).
edge(3304, 3305).
edge(3305, 3306).
edge(3306, 3307).
edge(3307, 3308).
edge(3308, 3309).
edge(3309, 3310).
edge(3310, 3311).
edge(3311, 3312).
edge(3312, 3313).
edge(3313, 3314).
edge(3314, 3315).
edge(3315, 3316).
edge(3316, 3317).
edge(3317, 3318).
edge(3318, 3319).
edge(3319, 3320).
edge(3320, 3321).
edge(3321, 3322).
edge(3322, 3323).
edge(3323, 3324).
edge(3324, 3325).
edge(3325, 3326).
edge(3326, 3327).
edge(3327, 3328).
edge(3328, 3329).
edge(3329, 3330).
edge(3330, 3331).
edge(3331, 3332).
edge(3332, 3333).
edge(3333, 3334).
edge(3334, 3335).
edge(3335, 3336).
edge(3336, 3337).
edge(3337, 3338).
edge(3338, 3339).
edge(3339, 3340).
edge(3340, 3341).
edge(3341, 3342).
edge(3342, 3343).
edge(3343, 3344).
edge(3344, 3345).
edge(3345, 3346).
edge(3346, 3347).
edge(3347, 3348).
edge(3348, 3349).
edge(3349, 3350).
edge(3350, 3351).
edge(3351, 3352).
edge(3352, 3353).
edge(3353, 3354).
edge(3354, 3355).
edge(3355, 3356).
edge(3356, 3357).
edge(3357, 3358).
edge(3358, 3359).
edge(3359, 3360).
edge(3360, 3361).
edge(3361, 3362).
edge(3362, 3363).
edge(3363, 3364).
edge(3364, 3365).
edge(3365, 3366).
edge(3366, 3367).
edge(3367, 3368).
edge(3368, 3369).
edge(3369, 3370).
edge(3370, 3371).
edge(3371, 3372).
edge(3372, 3373).
edge(3373, 3374).
edge(3374, 3375).
edge(3375, 3376).
edge(3376, 3377).
edge(3377, 3378).
edge(3378, 3379).
edge(3379, 3380).
edge(3380, 3381).
edge(3381, 3382).
edge(3382, 3383).
edge(3383, 3384).
edge(3384, 3385).
edge(3385, 3386).
edge(3386, 3387).
edge(3387, 3388).
edge(3388, 3389).
edge(3389, 3390).
edge(3390, 3391).
edge(3391, 3392).
edge(3392, 3393).
edge(3393, 3394).
edge(3394, 3395).
edge(3395, 3396).
edge(3396, 3397).
edge(3397, 3398).
edge(3398, 3399).
edge(3399, 3400).
edge(3400, 3401).
edge(3401, 3402).
edge(3402, 3403).
edge(3403, 3404).
edge(3404, 3405).
edge(3405, 3406).
edge(3406, 3407).
edge(3407, 3408).
edge(3408, 3409).
edge(3409, 3410).
edge(3410, 3411).
edge(3411, 3412).
edge(3412, 3413).
edge(3413, 3414).
edge(3414, 3415).
edge(3415, 3416).
edge(3416, 3417).
edge(3417, 3418).
edge(3418, 3419).
edge(3419, 3420).
edge(3420, 3421).
edge(3421, 3422).
edge(3422, 3423).
edge(3423, 3424).
edge(3424, 3425).
edge(3425, 3426).
edge(3426, 3427).
edge(3427, 3428).
edge(3428, 3429).
edge(3429, 3430).
edge(3430, 3431).
edge(3431, 3432).
edge(3432, 3433).
edge(3433, 3434).
edge(3434, 3435).
edge(3435, 3436).
edge(3436, 3437).
edge(3437, 3438).
edge(3438, 3439).
edge(3439, 3440).
edge(3440, 3441).
edge(3441, 3442).
edge(3442, 3443).
edge(3443, 3444).
edge(3444, 3445).
edge(3445, 3446).
edge(3446, 3447).
edge(3447, 3448).
edge(3448, 3449).
edge(3449, 3450).
edge(3450, 3451).
edge(3451, 3452).
edge(3452, 3453).
edge(3453, 3454).
edge(3454, 3455).
edge(3455, 3456).
edge(3456, 3457).
edge(3457, 3458).
edge(3458, 3459).
edge(3459, 3460).
edge(3460, 3461).
edge(3461, 3462).
edge(3462, 3463).
edge(3463, 3464).
edge(3464, 3465).
edge(3465, 3466).
edge(3466, 3467).
edge(3467, 3468).
edge(3468, 3469).
edge(3469, 3470).
edge(3470, 3471).
edge(3471, 3472).
edge(3472, 3473).
edge(3473, 3474).
edge(3474, 3475).
edge(3475, 3476).
edge(3476, 3477).
edge(3477, 3478).
edge(3478, 3479).
edge(3479, 3480).
edge(3480, 3481).
edge(3481, 3482).
edge(3482, 3483).
edge(3483, 3484).
edge(3484, 3485).
edge(3485, 3486).
edge(3486, 3487).
edge(3487, 3488).
edge(3488, 3489).
edge(3489, 3490).
edge(3490, 3491).
edge(3491, 3492).
edge(3492, 3493).
edge(3493, 3494).
edge(3494, 3495).
edge(3495, 3496).
edge(3496, 3497).
edge(3497, 3498).
edge(3498, 3499).
edge(3499, 3500).
edge(3500, 3501).
edge(3501, 3502).
edge(3502, 3503).
edge(3503, 3504).
edge(3504, 3505).
edge(3505, 3506).
edge(3506, 3507).
edge(3507, 3508).
edge(3508, 3509).
edge(3509, 3510).
edge(3510, 3511).
edge(3511, 3512).
edge(3512, 3513).
edge(3513, 3514).
edge(3514, 3515).
edge(3515, 3516).
edge(3516, 3517).
edge(3517, 3518).
edge(3518, 3519).
edge(3519, 3520).
edge(3520, 3521).
edge(3521, 3522).
edge(3522, 3523).
edge(3523, 3524).
edge(3524, 3525).
edge(3525, 3526).
edge(3526, 3527).
edge(3527, 3528).
edge(3528, 3529).
edge(3529, 3530).
edge(3530, 3531).
edge(3531, 3532).
edge(3532, 3533).
edge(3533, 3534).
edge(3534, 3535).
edge(3535, 3536).
edge(3536, 3537).
edge(3537, 3538).
edge(3538, 3539).
edge(3539, 3540).
edge(3540, 3541).
edge(3541, 3542).
edge(3542, 3543).
edge(3543, 3544).
edge(3544, 3545).
edge(3545, 3546).
edge(3546, 3547).
edge(3547, 3548).
edge(3548, 3549).
edge(3549, 3550).
edge(3550, 3551).
edge(3551, 3552).
edge(3552, 3553).
edge(3553, 3554).
edge(3554, 3555).
edge(3555, 3556).
edge(3556, 3557).
edge(3557, 3558).
edge(3558, 3559).
edge(3559, 3560).
edge(3560, 3561).
edge(3561, 3562).
edge(3562, 3563).
edge(3563, 3564).
edge(3564, 3565).
edge(3565, 3566).
edge(3566, 3567).
edge(3567, 3568).
edge(3568, 3569).
edge(3569, 3570).
edge(3570, 3571).
edge(3571, 3572).
edge(3572, 3573).
edge(3573, 3574).
edge(3574, 3575).
edge(3575, 3576).
edge(3576, 3577).
edge(3577, 3578).
edge(3578, 3579).
edge(3579, 3580).
edge(3580, 3581).
edge(3581, 3582).
edge(3582, 3583).
edge(3583, 3584).
edge(3584, 3585).
edge(3585, 3586).
edge(3586, 3587).
edge(3587, 3588).
edge(3588, 3589).
edge(3589, 3590).
edge(3590, 3591).
edge(3591, 3592).
edge(3592, 3593).
edge(3593, 3594).
edge(3594, 3595).
edge(3595, 3596).
edge(3596, 3597).
edge(3597, 3598).
edge(3598, 3599).
edge(3599, 3600).
edge(3600, 3601).
edge(3601, 3602).
edge(3602, 3603).
edge(3603, 3604).
edge(3604, 3605).
edge(3605, 3606).
edge(3606, 3607).
edge(3607, 3608).
edge(3608, 3609).
edge(3609, 3610).
edge(3610, 3611).
edge(3611, 3612).
edge(3612, 3613).
edge(3613, 3614).
edge(3614, 3615).
edge(3615, 3616).
edge(3616, 3617).
edge(3617, 3618).
edge(3618, 3619).
edge(3619, 3620).
edge(3620, 3621).
edge(3621, 3622).
edge(3622, 3623).
edge(3623, 3624).
edge(3624, 3625).
edge(3625, 3626).
edge(3626, 3627).
edge(3627, 3628).
edge(3628, 3629).
edge(3629, 3630).
edge(3630, 3631).
edge(3631, 3632).
edge(3632, 3633).
edge(3633, 3634).
edge(3634, 3635).
edge(3635, 3636).
edge(3636, 3637).
edge(3637, 3638).
edge(3638, 3639).
edge(3639, 3640).
edge(3640, 3641).
edge(3641, 3642).
edge(3642, 3643).
edge(3643, 3644).
edge(3644, 3645).
edge(3645, 3646).
edge(3646, 3647).
edge(3647, 3648).
edge(3648, 3649).
edge(3649, 3650).
edge(3650, 3651).
edge(3651, 3652).
edge(3652, 3653).
edge(3653, 3654).
edge(3654, 3655).
edge(3655, 3656).
edge(3656, 3657).
edge(3657, 3658).
edge(3658, 3659).
edge(3659, 3660).
edge(3660, 3661).
edge(3661, 3662).
edge(3662, 3663).
edge(3663, 3664).
edge(3664, 3665).
edge(3665, 3666).
edge(3666, 3667).
edge(3667, 3668).
edge(3668, 3669).
edge(3669, 3670).
edge(3670, 3671).
edge(3671, 3672).
edge(3672, 3673).
edge(3673, 3674).
edge(3674, 3675).
edge(3675, 3676).
edge(3676, 3677).
edge(3677, 3678).
edge(3678, 3679).
edge(3679, 3680).
edge(3680, 3681).
edge(3681, 3682).
edge(3682, 3683).
edge(3683, 3684).
edge(3684, 3685).
edge(3685, 3686).
edge(3686, 3687).
edge(3687, 3688).
edge(3688, 3689).
edge(3689, 3690).
edge(3690, 3691).
edge(3691, 3692).
edge(3692, 3693).
edge(3693, 3694).
edge(3694, 3695).
edge(3695, 3696).
edge(3696, 3697).
edge(3697, 3698).
edge(3698, 3699).
edge(3699, 3700).
edge(3700, 3701).
edge(3701, 3702).
edge(3702, 3703).
edge(3703, 3704).
edge(3704, 3705).
edge(3705, 3706).
edge(3706, 3707).
edge(3707, 3708).
edge(3708, 3709).
edge(3709, 3710).
edge(3710, 3711).
edge(3711, 3712).
edge(3712, 3713).
edge(3713, 3714).
edge(3714, 3715).
edge(3715, 3716).
edge(3716, 3717).
edge(3717, 3718).
edge(3718, 3719).
edge(3719, 3720).
edge(3720, 3721).
edge(3721, 3722).
edge(3722, 3723).
edge(3723, 3724).
edge(3724, 3725).
edge(3725, 3726).
edge(3726, 3727).
edge(3727, 3728).
edge(3728, 3729).
edge(3729, 3730).
edge(3730, 3731).
edge(3731, 3732).
edge(3732, 3733).
edge(3733, 3734).
edge(3734, 3735).
edge(3735, 3736).
edge(3736, 3737).
edge(3737, 3738).
edge(3738, 3739).
edge(3739, 3740).
edge(3740, 3741).
edge(3741, 3742).
edge(3742, 3743).
edge(3743, 3744).
edge(3744, 3745).
edge(3745, 3746).
edge(3746, 3747).
edge(3747, 3748).
edge(3748, 3749).
edge(3749, 3750).
edge(3750, 3751).
edge(3751, 3752).
edge(3752, 3753).
edge(3753, 3754).
edge(3754, 3755).
edge(3755, 3756).
edge(3756, 3757).
edge(3757, 3758).
edge(3758, 3759).
edge(3759, 3760).
edge(3760, 3761).
edge(3761, 3762).
edge(3762, 3763).
edge(3763, 3764).
edge(3764, 3765).
edge(3765, 3766).
edge(3766, 3767).
edge(3767, 3768).
edge(3768, 3769).
edge(3769, 3770).
edge(3770, 3771).
edge(3771, 3772).
edge(3772, 3773).
edge(3773, 3774).
edge(3774, 3775).
edge(3775, 3776).
edge(3776, 3777).
edge(3777, 3778).
edge(3778, 3779).
edge(3779, 3780).
edge(3780, 3781).
edge(3781, 3782).
edge(3782, 3783).
edge(3783, 3784).
edge(3784, 3785).
edge(3785, 3786).
edge(3786, 3787).
edge(3787, 3788).
edge(3788, 3789).
edge(3789, 3790).
edge(3790, 3791).
edge(3791, 3792).
edge(3792, 3793).
edge(3793, 3794).
edge(3794, 3795).
edge(3795, 3796).
edge(3796, 3797).
edge(3797, 3798).
edge(3798, 3799).
edge(3799, 3800).
edge(3800, 3801).
edge(3801, 3802).
edge(3802, 3803).
edge(3803, 3804).
edge(3804, 3805).
edge(3805, 3806).
edge(3806, 3807).
edge(3807, 3808).
edge(3808, 3809).
edge(3809, 3810).
edge(3810, 3811).
edge(3811, 3812).
edge(3812, 3813).
edge(3813, 3814).
edge(3814, 3815).
edge(3815, 3816).
edge(3816, 3817).
edge(3817, 3818).
edge(3818, 3819).
edge(3819, 3820).
edge(3820, 3821).
edge(3821, 3822).
edge(3822, 3823).
edge(3823, 3824).
edge(3824, 3825).
edge(3825, 3826).
edge(3826, 3827).
edge(3827, 3828).
edge(3828, 3829).
edge(3829, 3830).
edge(3830, 3831).
edge(3831, 3832).
edge(3832, 3833).
edge(3833, 3834).
edge(3834, 3835).
edge(3835, 3836).
edge(3836, 3837).
edge(3837, 3838).
edge(3838, 3839).
edge(3839, 3840).
edge(3840, 3841).
edge(3841, 3842).
edge(3842, 3843).
edge(3843, 3844).
edge(3844, 3845).
edge(3845, 3846).
edge(3846, 3847).
edge(3847, 3848).
edge(3848, 3849).
edge(3849, 3850).
edge(3850, 3851).
edge(3851, 3852).
edge(3852, 3853).
edge(3853, 3854).
edge(3854, 3855).
edge(3855, 3856).
edge(3856, 3857).
edge(3857, 3858).
edge(3858, 3859).
edge(3859, 3860).
edge(3860, 3861).
edge(3861, 3862).
edge(3862, 3863).
edge(3863, 3864).
edge(3864, 3865).
edge(3865, 3866).
edge(3866, 3867).
edge(3867, 3868).
edge(3868, 3869).
edge(3869, 3870).
edge(3870, 3871).
edge(3871, 3872).
edge(3872, 3873).
edge(3873, 3874).
edge(3874, 3875).
edge(3875, 3876).
edge(3876, 3877).
edge(3877, 3878).
edge(3878, 3879).
edge(3879, 3880).
edge(3880, 3881).
edge(3881, 3882).
edge(3882, 3883).
edge(3883, 3884).
edge(3884, 3885).
edge(3885, 3886).
edge(3886, 3887).
edge(3887, 3888).
edge(3888, 3889).
edge(3889, 3890).
edge(3890, 3891).
edge(3891, 3892).
edge(3892, 3893).
edge(3893, 3894).
edge(3894, 3895).
edge(3895, 3896).
edge(3896, 3897).
edge(3897, 3898).
edge(3898, 3899).
edge(3899, 3900).
edge(3900, 3901).
edge(3901, 3902).
edge(3902, 3903).
edge(3903, 3904).
edge(3904, 3905).
edge(3905, 3906).
edge(3906, 3907).
edge(3907, 3908).
edge(3908, 3909).
edge(3909, 3910).
edge(3910, 3911).
edge(3911, 3912).
edge(3912, 3913).
edge(3913, 3914).
edge(3914, 3915).
edge(3915, 3916).
edge(3916, 3917).
edge(3917, 3918).
edge(3918, 3919).
edge(3919, 3920).
edge(3920, 3921).
edge(3921, 3922).
edge(3922, 3923).
edge(3923, 3924).
edge(3924, 3925).
edge(3925, 3926).
edge(3926, 3927).
edge(3927, 3928).
edge(3928, 3929).
edge(3929, 3930).
edge(3930, 3931).
edge(3931, 3932).
edge(3932, 3933).
edge(3933, 3934).
edge(3934, 3935).
edge(3935, 3936).
edge(3936, 3937).
edge(3937, 3938).
edge(3938, 3939).
edge(3939, 3940).
edge(3940, 3941).
edge(3941, 3942).
edge(3942, 3943).
edge(3943, 3944).
edge(3944, 3945).
edge(3945, 3946).
edge(3946, 3947).
edge(3947, 3948).
edge(3948, 3949).
edge(3949, 3950).
edge(3950, 3951).
edge(3951, 3952).
edge(3952, 3953).
edge(3953, 3954).
edge(3954, 3955).
edge(3955, 3956).
edge(3956, 3957).
edge(3957, 3958).
edge(3958, 3959).
edge(3959, 3960).
edge(3960, 3961).
edge(3961, 3962).
edge(3962, 3963).
edge(3963, 3964).
edge(3964, 3965).
edge(3965, 3966).
edge(3966, 3967).
edge(3967, 3968).
edge(3968, 3969).
edge(3969, 3970).
edge(3970, 3971).
edge(3971, 3972).
edge(3972, 3973).
edge(3973, 3974).
edge(3974, 3975).
edge(3975, 3976).
edge(3976, 3977).
edge(3977, 3978).
edge(3978, 3979).
edge(3979, 3980).
edge(3980, 3981).
edge(3981, 3982).
edge(3982, 3983).
edge(3983, 3984).
edge(3984, 3985).
edge(3985, 3986).
edge(3986, 3987).
edge(3987, 3988).
edge(3988, 3989).
edge(3989, 3990).
edge(3990, 3991).
edge(3991, 3992).
edge(3992, 3993).
edge(3993, 3994).
edge(3994, 3995).
edge(3995, 3996).
edge(3996, 3997).
edge(3997, 3998).
edge(3998, 3999).
edge(3999, 4000).
edge(4000, 4001).
edge(4001, 4002).
edge(4002, 4003).
edge(4003, 4004).
edge(4004, 4005).
edge(4005, 4006).
edge(4006, 4007).
edge(4007, 4008).
edge(4008, 4009).
edge(4009, 4010).
edge(4010, 4011).
edge(4011, 4012).
edge(4012, 4013).
edge(4013, 4014).
edge(4014, 4015).
edge(4015, 4016).
edge(4016, 4017).
edge(4017, 4018).
edge(4018, 4019).
edge(4019, 4020).
edge(4020, 4021).
edge(4021, 4022).
edge(4022, 4023).
edge(4023, 4024).
edge(4024, 4025).
edge(4025, 4026).
edge(4026, 4027).
edge(4027, 4028).
edge(4028, 4029).
edge(4029, 4030).
edge(4030, 4031).
edge(4031, 4032).
edge(4032, 4033).
edge(4033, 4034).
edge(4034, 4035).
edge(4035, 4036).
edge(4036, 4037).
edge(4037, 4038).
edge(4038, 4039).
edge(4039, 4040).
edge(4040, 4041).
edge(4041, 4042).
edge(4042, 4043).
edge(4043, 4044).
edge(4044, 4045).
edge(4045, 4046).
edge(4046, 4047).
edge(4047, 4048).
edge(4048, 4049).
edge(4049, 4050).
edge(4050, 4051).
edge(4051, 4052).
edge(4052, 4053).
edge(4053, 4054).
edge(4054, 4055).
edge(4055, 4056).
edge(4056, 4057).
edge(4057, 4058).
edge(4058, 4059).
edge(4059, 4060).
edge(4060, 4061).
edge(4061, 4062).
edge(4062, 4063).
edge(4063, 4064).
edge(4064, 4065).
edge(4065, 4066).
edge(4066, 4067).
edge(4067, 4068).
edge(4068, 4069).
edge(4069, 4070).
edge(4070, 4071).
edge(4071, 4072).
edge(4072, 4073).
edge(4073, 4074).
edge(4074, 4075).
edge(4075, 4076).
edge(4076, 4077).
edge(4077, 4078).
edge(4078, 4079).
edge(4079, 4080).
edge(4080, 4081).
edge(4081, 4082).
edge(4082, 4083).
edge(4083, 4084).
edge(4084, 4085).
edge(4085, 4086).
edge(4086, 4087).
edge(4087, 4088).
edge(4088, 4089).
edge(4089, 4090).
edge(4090, 4091).
edge(4091, 4092).
edge(4092, 4093).
edge(4093, 4094).
edge(4094, 4095).
edge(4095, 4096).
edge(4096, 4097).
edge(4097, 4098).
edge(4098, 4099).
edge(4099, 4100).
edge(4100, 4101).
edge(4101, 4102).
edge(4102, 4103).
edge(4103, 4104).
edge(4104, 4105).
edge(4105, 4106).
edge(4106, 4107).
edge(4107, 4108).
edge(4108, 4109).
edge(4109, 4110).
edge(4110, 4111).
edge(4111, 4112).
edge(4112, 4113).
edge(4113, 4114).
edge(4114, 4115).
edge(4115, 4116).
edge(4116, 4117).
edge(4117, 4118).
edge(4118, 4119).
edge(4119, 4120).
edge(4120, 4121).
edge(4121, 4122).
edge(4122, 4123).
edge(4123, 4124).
edge(4124, 4125).
edge(4125, 4126).
edge(4126, 4127).
edge(4127, 4128).
edge(4128, 4129).
edge(4129, 4130).
edge(4130, 4131).
edge(4131, 4132).
edge(4132, 4133).
edge(4133, 4134).
edge(4134, 4135).
edge(4135, 4136).
edge(4136, 4137).
edge(4137, 4138).
edge(4138, 4139).
edge(4139, 4140).
edge(4140, 4141).
edge(4141, 4142).
edge(4142, 4143).
edge(4143, 4144).
edge(4144, 4145).
edge(4145, 4146).
edge(4146, 4147).
edge(4147, 4148).
edge(4148, 4149).
edge(4149, 4150).
edge(4150, 4151).
edge(4151, 4152).
edge(4152, 4153).
edge(4153, 4154).
edge(4154, 4155).
edge(4155, 4156).
edge(4156, 4157).
edge(4157, 4158).
edge(4158, 4159).
edge(4159, 4160).
edge(4160, 4161).
edge(4161, 4162).
edge(4162, 4163).
edge(4163, 4164).
edge(4164, 4165).
edge(4165, 4166).
edge(4166, 4167).
edge(4167, 4168).
edge(4168, 4169).
edge(4169, 4170).
edge(4170, 4171).
edge(4171, 4172).
edge(4172, 4173).
edge(4173, 4174).
edge(4174, 4175).
edge(4175, 4176).
edge(4176, 4177).
edge(4177, 4178).
edge(4178, 4179).
edge(4179, 4180).
edge(4180, 4181).
edge(4181, 4182).
edge(4182, 4183).
edge(4183, 4184).
edge(4184, 4185).
edge(4185, 4186).
edge(4186, 4187).
edge(4187, 4188).
edge(4188, 4189).
edge(4189, 4190).
edge(4190, 4191).
edge(4191, 4192).
edge(4192, 4193).
edge(4193, 4194).
edge(4194, 4195).
edge(4195, 4196).
edge(4196, 4197).
edge(4197, 4198).
edge(4198, 4199).
edge(4199, 4200).
edge(4200, 4201).
edge(4201, 4202).
edge(4202, 4203).
edge(4203, 4204).
edge(4204, 4205).
edge(4205, 4206).
edge(4206, 4207).
edge(4207, 4208).
edge(4208, 4209).
edge(4209, 4210).
edge(4210, 4211).
edge(4211, 4212).
edge(4212, 4213).
edge(4213, 4214).
edge(4214, 4215).
edge(4215, 4216).
edge(4216, 4217).
edge(4217, 4218).
edge(4218, 4219).
edge(4219, 4220).
edge(4220, 4221).
edge(4221, 4222).
edge(4222, 4223).
edge(4223, 4224).
edge(4224, 4225).
edge(4225, 4226).
edge(4226, 4227).
edge(4227, 4228).
edge(4228, 4229).
edge(4229, 4230).
edge(4230, 4231).
edge(4231, 4232).
edge(4232, 4233).
edge(4233, 4234).
edge(4234, 4235).
edge(4235, 4236).
edge(4236, 4237).
edge(4237, 4238).
edge(4238, 4239).
edge(4239, 4240).
edge(4240, 4241).
edge(4241, 4242).
edge(4242, 4243).
edge(4243, 4244).
edge(4244, 4245).
edge(4245, 4246).
edge(4246, 4247).
edge(4247, 4248).
edge(4248, 4249).
edge(4249, 4250).
edge(4250, 4251).
edge(4251, 4252).
edge(4252, 4253).
edge(4253, 4254).
edge(4254, 4255).
edge(4255, 4256).
edge(4256, 4257).
edge(4257, 4258).
edge(4258, 4259).
edge(4259, 4260).
edge(4260, 4261).
edge(4261, 4262).
edge(4262, 4263).
edge(4263, 4264).
edge(4264, 4265).
edge(4265, 4266).
edge(4266, 4267).
edge(4267, 4268).
edge(4268, 4269).
edge(4269, 4270).
edge(4270, 4271).
edge(4271, 4272).
edge(4272, 4273).
edge(4273, 4274).
edge(4274, 4275).
edge(4275, 4276).
edge(4276, 4277).
edge(4277, 4278).
edge(4278, 4279).
edge(4279, 4280).
edge(4280, 4281).
edge(4281, 4282).
edge(4282, 4283).
edge(4283, 4284).
edge(4284, 4285).
edge(4285, 4286).
edge(4286, 4287).
edge(4287, 4288).
edge(4288, 4289).
edge(4289, 4290).
edge(4290, 4291).
edge(4291, 4292).
edge(4292, 4293).
edge(4293, 4294).
edge(4294, 4295).
edge(4295, 4296).
edge(4296, 4297).
edge(4297, 4298).
edge(4298, 4299).
edge(4299, 4300).
edge(4300, 4301).
edge(4301, 4302).
edge(4302, 4303).
edge(4303, 4304).
edge(4304, 4305).
edge(4305, 4306).
edge(4306, 4307).
edge(4307, 4308).
edge(4308, 4309).
edge(4309, 4310).
edge(4310, 4311).
edge(4311, 4312).
edge(4312, 4313).
edge(4313, 4314).
edge(4314, 4315).
edge(4315, 4316).
edge(4316, 4317).
edge(4317, 4318).
edge(4318, 4319).
edge(4319, 4320).
edge(4320, 4321).
edge(4321, 4322).
edge(4322, 4323).
edge(4323, 4324).
edge(4324, 4325).
edge(4325, 4326).
edge(4326, 4327).
edge(4327, 4328).
edge(4328, 4329).
edge(4329, 4330).
edge(4330, 4331).
edge(4331, 4332).
edge(4332, 4333).
edge(4333, 4334).
edge(4334, 4335).
edge(4335, 4336).
edge(4336, 4337).
edge(4337, 4338).
edge(4338, 4339).
edge(4339, 4340).
edge(4340, 4341).
edge(4341, 4342).
edge(4342, 4343).
edge(4343, 4344).
edge(4344, 4345).
edge(4345, 4346).
edge(4346, 4347).
edge(4347, 4348).
edge(4348, 4349).
edge(4349, 4350).
edge(4350, 4351).
edge(4351, 4352).
edge(4352, 4353).
edge(4353, 4354).
edge(4354, 4355).
edge(4355, 4356).
edge(4356, 4357).
edge(4357, 4358).
edge(4358, 4359).
edge(4359, 4360).
edge(4360, 4361).
edge(4361, 4362).
edge(4362, 4363).
edge(4363, 4364).
edge(4364, 4365).
edge(4365, 4366).
edge(4366, 4367).
edge(4367, 4368).
edge(4368, 4369).
edge(4369, 4370).
edge(4370, 4371).
edge(4371, 4372).
edge(4372, 4373).
edge(4373, 4374).
edge(4374, 4375).
edge(4375, 4376).
edge(4376, 4377).
edge(4377, 4378).
edge(4378, 4379).
edge(4379, 4380).
edge(4380, 4381).
edge(4381, 4382).
edge(4382, 4383).
edge(4383, 4384).
edge(4384, 4385).
edge(4385, 4386).
edge(4386, 4387).
edge(4387, 4388).
edge(4388, 4389).
edge(4389, 4390).
edge(4390, 4391).
edge(4391, 4392).
edge(4392, 4393).
edge(4393, 4394).
edge(4394, 4395).
edge(4395, 4396).
edge(4396, 4397).
edge(4397, 4398).
edge(4398, 4399).
edge(4399, 4400).
edge(4400, 4401).
edge(4401, 4402).
edge(4402, 4403).
edge(4403, 4404).
edge(4404, 4405).
edge(4405, 4406).
edge(4406, 4407).
edge(4407, 4408).
edge(4408, 4409).
edge(4409, 4410).
edge(4410, 4411).
edge(4411, 4412).
edge(4412, 4413).
edge(4413, 4414).
edge(4414, 4415).
edge(4415, 4416).
edge(4416, 4417).
edge(4417, 4418).
edge(4418, 4419).
edge(4419, 4420).
edge(4420, 4421).
edge(4421, 4422).
edge(4422, 4423).
edge(4423, 4424).
edge(4424, 4425).
edge(4425, 4426).
edge(4426, 4427).
edge(4427, 4428).
edge(4428, 4429).
edge(4429, 4430).
edge(4430, 4431).
edge(4431, 4432).
edge(4432, 4433).
edge(4433, 4434).
edge(4434, 4435).
edge(4435, 4436).
edge(4436, 4437).
edge(4437, 4438).
edge(4438, 4439).
edge(4439, 4440).
edge(4440, 4441).
edge(4441, 4442).
edge(4442, 4443).
edge(4443, 4444).
edge(4444, 4445).
edge(4445, 4446).
edge(4446, 4447).
edge(4447, 4448).
edge(4448, 4449).
edge(4449, 4450).
edge(4450, 4451).
edge(4451, 4452).
edge(4452, 4453).
edge(4453, 4454).
edge(4454, 4455).
edge(4455, 4456).
edge(4456, 4457).
edge(4457, 4458).
edge(4458, 4459).
edge(4459, 4460).
edge(4460, 4461).
edge(4461, 4462).
edge(4462, 4463).
edge(4463, 4464).
edge(4464, 4465).
edge(4465, 4466).
edge(4466, 4467).
edge(4467, 4468).
edge(4468, 4469).
edge(4469, 4470).
edge(4470, 4471).
edge(4471, 4472).
edge(4472, 4473).
edge(4473, 4474).
edge(4474, 4475).
edge(4475, 4476).
edge(4476, 4477).
edge(4477, 4478).
edge(4478, 4479).
edge(4479, 4480).
edge(4480, 4481).
edge(4481, 4482).
edge(4482, 4483).
edge(4483, 4484).
edge(4484, 4485).
edge(4485, 4486).
edge(4486, 4487).
edge(4487, 4488).
edge(4488, 4489).
edge(4489, 4490).
edge(4490, 4491).
edge(4491, 4492).
edge(4492, 4493).
edge(4493, 4494).
edge(4494, 4495).
edge(4495, 4496).
edge(4496, 4497).
edge(4497, 4498).
edge(4498, 4499).
edge(4499, 4500).
edge(4500, 4501).
edge(4501, 4502).
edge(4502, 4503).
edge(4503, 4504).
edge(4504, 4505).
edge(4505, 4506).
edge(4506, 4507).
edge(4507, 4508).
edge(4508, 4509).
edge(4509, 4510).
edge(4510, 4511).
edge(4511, 4512).
edge(4512, 4513).
edge(4513, 4514).
edge(4514, 4515).
edge(4515, 4516).
edge(4516, 4517).
edge(4517, 4518).
edge(4518, 4519).
edge(4519, 4520).
edge(4520, 4521).
edge(4521, 4522).
edge(4522, 4523).
edge(4523, 4524).
edge(4524, 4525).
edge(4525, 4526).
edge(4526, 4527).
edge(4527, 4528).
edge(4528, 4529).
edge(4529, 4530).
edge(4530, 4531).
edge(4531, 4532).
edge(4532, 4533).
edge(4533, 4534).
edge(4534, 4535).
edge(4535, 4536).
edge(4536, 4537).
edge(4537, 4538).
edge(4538, 4539).
edge(4539, 4540).
edge(4540, 4541).
edge(4541, 4542).
edge(4542, 4543).
edge(4543, 4544).
edge(4544, 4545).
edge(4545, 4546).
edge(4546, 4547).
edge(4547, 4548).
edge(4548, 4549).
edge(4549, 4550).
edge(4550, 4551).
edge(4551, 4552).
edge(4552, 4553).
edge(4553, 4554).
edge(4554, 4555).
edge(4555, 4556).
edge(4556, 4557).
edge(4557, 4558).
edge(4558, 4559).
edge(4559, 4560).
edge(4560, 4561).
edge(4561, 4562).
edge(4562, 4563).
edge(4563, 4564).
edge(4564, 4565).
edge(4565, 4566).
edge(4566, 4567).
edge(4567, 4568).
edge(4568, 4569).
edge(4569, 4570).
edge(4570, 4571).
edge(4571, 4572).
edge(4572, 4573).
edge(4573, 4574).
edge(4574, 4575).
edge(4575, 4576).
edge(4576, 4577).
edge(4577, 4578).
edge(4578, 4579).
edge(4579, 4580).
edge(4580, 4581).
edge(4581, 4582).
edge(4582, 4583).
edge(4583, 4584).
edge(4584, 4585).
edge(4585, 4586).
edge(4586, 4587).
edge(4587, 4588).
edge(4588, 4589).
edge(4589, 4590).
edge(4590, 4591).
edge(4591, 4592).
edge(4592, 4593).
edge(4593, 4594).
edge(4594, 4595).
edge(4595, 4596).
edge(4596, 4597).
edge(4597, 4598).
edge(4598, 4599).
edge(4599, 4600).
edge(4600, 4601).
edge(4601, 4602).
edge(4602, 4603).
edge(4603, 4604).
edge(4604, 4605).
edge(4605, 4606).
edge(4606, 4607).
edge(4607, 4608).
edge(4608, 4609).
edge(4609, 4610).
edge(4610, 4611).
edge(4611, 4612).
edge(4612, 4613).
edge(4613, 4614).
edge(4614, 4615).
edge(4615, 4616).
edge(4616, 4617).
edge(4617, 4618).
edge(4618, 4619).
edge(4619, 4620).
edge(4620, 4621).
edge(4621, 4622).
edge(4622, 4623).
edge(4623, 4624).
edge(4624, 4625).
edge(4625, 4626).
edge(4626, 4627).
edge(4627, 4628).
edge(4628, 4629).
edge(4629, 4630).
edge(4630, 4631).
edge(4631, 4632).
edge(4632, 4633).
edge(4633, 4634).
edge(4634, 4635).
edge(4635, 4636).
edge(4636, 4637).
edge(4637, 4638).
edge(4638, 4639).
edge(4639, 4640).
edge(4640, 4641).
edge(4641, 4642).
edge(4642, 4643).
edge(4643, 4644).
edge(4644, 4645).
edge(4645, 4646).
edge(4646, 4647).
edge(4647, 4648).
edge(4648, 4649).
edge(4649, 4650).
edge(4650, 4651).
edge(4651, 4652).
edge(4652, 4653).
edge(4653, 4654).
edge(4654, 4655).
edge(4655, 4656).
edge(4656, 4657).
edge(4657, 4658).
edge(4658, 4659).
edge(4659, 4660).
edge(4660, 4661).
edge(4661, 4662).
edge(4662, 4663).
edge(4663, 4664).
edge(4664, 4665).
edge(4665, 4666).
edge(4666, 4667).
edge(4667, 4668).
edge(4668, 4669).
edge(4669, 4670).
edge(4670, 4671).
edge(4671, 4672).
edge(4672, 4673).
edge(4673, 4674).
edge(4674, 4675).
edge(4675, 4676).
edge(4676, 4677).
edge(4677, 4678).
edge(4678, 4679).
edge(4679, 4680).
edge(4680, 4681).
edge(4681, 4682).
edge(4682, 4683).
edge(4683, 4684).
edge(4684, 4685).
edge(4685, 4686).
edge(4686, 4687).
edge(4687, 4688).
edge(4688, 4689).
edge(4689, 4690).
edge(4690, 4691).
edge(4691, 4692).
edge(4692, 4693).
edge(4693, 4694).
edge(4694, 4695).
edge(4695, 4696).
edge(4696, 4697).
edge(4697, 4698).
edge(4698, 4699).
edge(4699, 4700).
edge(4700, 4701).
edge(4701, 4702).
edge(4702, 4703).
edge(4703, 4704).
edge(4704, 4705).
edge(4705, 4706).
edge(4706, 4707).
edge(4707, 4708).
edge(4708, 4709).
edge(4709, 4710).
edge(4710, 4711).
edge(4711, 4712).
edge(4712, 4713).
edge(4713, 4714).
edge(4714, 4715).
edge(4715, 4716).
edge(4716, 4717).
edge(4717, 4718).
edge(4718, 4719).
edge(4719, 4720).
edge(4720, 4721).
edge(4721, 4722).
edge(4722, 4723).
edge(4723, 4724).
edge(4724, 4725).
edge(4725, 4726).
edge(4726, 4727).
edge(4727, 4728).
edge(4728, 4729).
edge(4729, 4730).
edge(4730, 4731).
edge(4731, 4732).
edge(4732, 4733).
edge(4733, 4734).
edge(4734, 4735).
edge(4735, 4736).
edge(4736, 4737).
edge(4737, 4738).
edge(4738, 4739).
edge(4739, 4740).
edge(4740, 4741).
edge(4741, 4742).
edge(4742, 4743).
edge(4743, 4744).
edge(4744, 4745).
edge(4745, 4746).
edge(4746, 4747).
edge(4747, 4748).
edge(4748, 4749).
edge(4749, 4750).
edge(4750, 4751).
edge(4751, 4752).
edge(4752, 4753).
edge(4753, 4754).
edge(4754, 4755).
edge(4755, 4756).
edge(4756, 4757).
edge(4757, 4758).
edge(4758, 4759).
edge(4759, 4760).
edge(4760, 4761).
edge(4761, 4762).
edge(4762, 4763).
edge(4763, 4764).
edge(4764, 4765).
edge(4765, 4766).
edge(4766, 4767).
edge(4767, 4768).
edge(4768, 4769).
edge(4769, 4770).
edge(4770, 4771).
edge(4771, 4772).
edge(4772, 4773).
edge(4773, 4774).
edge(4774, 4775).
edge(4775, 4776).
edge(4776, 4777).
edge(4777, 4778).
edge(4778, 4779).
edge(4779, 4780).
edge(4780, 4781).
edge(4781, 4782).
edge(4782, 4783).
edge(4783, 4784).
edge(4784, 4785).
edge(4785, 4786).
edge(4786, 4787).
edge(4787, 4788).
edge(4788, 4789).
edge(4789, 4790).
edge(4790, 4791).
edge(4791, 4792).
edge(4792, 4793).
edge(4793, 4794).
edge(4794, 4795).
edge(4795, 4796).
edge(4796, 4797).
edge(4797, 4798).
edge(4798, 4799).
edge(4799, 4800).
edge(4800, 4801).
edge(4801, 4802).
edge(4802, 4803).
edge(4803, 4804).
edge(4804, 4805).
edge(4805, 4806).
edge(4806, 4807).
edge(4807, 4808).
edge(4808, 4809).
edge(4809, 4810).
edge(4810, 4811).
edge(4811, 4812).
edge(4812, 4813).
edge(4813, 4814).
edge(4814, 4815).
edge(4815, 4816).
edge(4816, 4817).
edge(4817, 4818).
edge(4818, 4819).
edge(4819, 4820).
edge(4820, 4821).
edge(4821, 4822).
edge(4822, 4823).
edge(4823, 4824).
edge(4824, 4825).
edge(4825, 4826).
edge(4826, 4827).
edge(4827, 4828).
edge(4828, 4829).
edge(4829, 4830).
edge(4830, 4831).
edge(4831, 4832).
edge(4832, 4833).
edge(4833, 4834).
edge(4834, 4835).
edge(4835, 4836).
edge(4836, 4837).
edge(4837, 4838).
edge(4838, 4839).
edge(4839, 4840).
edge(4840, 4841).
edge(4841, 4842).
edge(4842, 4843).
edge(4843, 4844).
edge(4844, 4845).
edge(4845, 4846).
edge(4846, 4847).
edge(4847, 4848).
edge(4848, 4849).
edge(4849, 4850).
edge(4850, 4851).
edge(4851, 4852).
edge(4852, 4853).
edge(4853, 4854).
edge(4854, 4855).
edge(4855, 4856).
edge(4856, 4857).
edge(4857, 4858).
edge(4858, 4859).
edge(4859, 4860).
edge(4860, 4861).
edge(4861, 4862).
edge(4862, 4863).
edge(4863, 4864).
edge(4864, 4865).
edge(4865, 4866).
edge(4866, 4867).
edge(4867, 4868).
edge(4868, 4869).
edge(4869, 4870).
edge(4870, 4871).
edge(4871, 4872).
edge(4872, 4873).
edge(4873, 4874).
edge(4874, 4875).
edge(4875, 4876).
edge(4876, 4877).
edge(4877, 4878).
edge(4878, 4879).
edge(4879, 4880).
edge(4880, 4881).
edge(4881, 4882).
edge(4882, 4883).
edge(4883, 4884).
edge(4884, 4885).
edge(4885, 4886).
edge(4886, 4887).
edge(4887, 4888).
edge(4888, 4889).
edge(4889, 4890).
edge(4890, 4891).
edge(4891, 4892).
edge(4892, 4893).
edge(4893, 4894).
edge(4894, 4895).
edge(4895, 4896).
edge(4896, 4897).
edge(4897, 4898).
edge(4898, 4899).
edge(4899, 4900).
edge(4900, 4901).
edge(4901, 4902).
edge(4902, 4903).
edge(4903, 4904).
edge(4904, 4905).
edge(4905, 4906).
edge(4906, 4907).
edge(4907, 4908).
edge(4908, 4909).
edge(4909, 4910).
edge(4910, 4911).
edge(4911, 4912).
edge(4912, 4913).
edge(4913, 4914).
edge(4914, 4915).
edge(4915, 4916).
edge(4916, 4917).
edge(4917, 4918).
edge(4918, 4919).
edge(4919, 4920).
edge(4920, 4921).
edge(4921, 4922).
edge(4922, 4923).
edge(4923, 4924).
edge(4924, 4925).
edge(4925, 4926).
edge(4926, 4927).
edge(4927, 4928).
edge(4928, 4929).
edge(4929, 4930).
edge(4930, 4931).
edge(4931, 4932).
edge(4932, 4933).
edge(4933, 4934).
edge(4934, 4935).
edge(4935, 4936).
edge(4936, 4937).
edge(4937, 4938).
edge(4938, 4939).
edge(4939, 4940).
edge(4940, 4941).
edge(4941, 4942).
edge(4942, 4943).
edge(4943, 4944).
edge(4944, 4945).
edge(4945, 4946).
edge(4946, 4947).
edge(4947, 4948).
edge(4948, 4949).
edge(4949, 4950).
edge(4950, 4951).
edge(4951, 4952).
edge(4952, 4953).
edge(4953, 4954).
edge(4954, 4955).
edge(4955, 4956).
edge(4956, 4957).
edge(4957, 4958).
edge(4958, 4959).
edge(4959, 4960).
edge(4960, 4961).
edge(4961, 4962).
edge(4962, 4963).
edge(4963, 4964).
edge(4964, 4965).
edge(4965, 4966).
edge(4966, 4967).
edge(4967, 4968).
edge(4968, 4969).
edge(4969, 4970).
edge(4970, 4971).
edge(4971, 4972).
edge(4972, 4973).
edge(4973, 4974).
edge(4974, 4975).
edge(4975, 4976).
edge(4976, 4977).
edge(4977, 4978).
edge(4978, 4979).
edge(4979, 4980).
edge(4980, 4981).
edge(4981, 4982).
edge(4982, 4983).
edge(4983, 4984).
edge(4984, 4985).
edge(4985, 4986).
edge(4986, 4987).
edge(4987, 4988).
edge(4988, 4989).
edge(4989, 4990).
edge(4990, 4991).
edge(4991, 4992).
edge(4992, 4993).
edge(4993, 4994).
edge(4994, 4995).
edge(4995, 4996).
edge(4996, 4997).
edge(4997, 4998).
edge(4998, 4999).
edge(4999, 5000).
edge(5000, 5001).
edge(5001, 5002).
edge(5002, 5003).
edge(5003, 5004).
edge(5004, 5005).
edge(5005, 5006).
edge(5006, 5007).
edge(5007, 5008).
edge(5008, 5009).
edge(5009, 5010).
edge(5010, 5011).
edge(5011, 5012).
edge(5012, 5013).
edge(5013, 5014).
edge(5014, 5015).
edge(5015, 5016).
edge(5016, 5017).
edge(5017, 5018).
edge(5018, 5019).
edge(5019, 5020).
edge(5020, 5021).
edge(5021, 5022).
edge(5022, 5023).
edge(5023, 5024).
edge(5024, 5025).
edge(5025, 5026).
edge(5026, 5027).
edge(5027, 5028).
edge(5028, 5029).
edge(5029, 5030).
edge(5030, 5031).
edge(5031, 5032).
edge(5032, 5033).
edge(5033, 5034).
edge(5034, 5035).
edge(5035, 5036).
edge(5036, 5037).
edge(5037, 5038).
edge(5038, 5039).
edge(5039, 5040).
edge(5040, 5041).
edge(5041, 5042).
edge(5042, 5043).
edge(5043, 5044).
edge(5044, 5045).
edge(5045, 5046).
edge(5046, 5047).
edge(5047, 5048).
edge(5048, 5049).
edge(5049, 5050).
edge(5050, 5051).
edge(5051, 5052).
edge(5052, 5053).
edge(5053, 5054).
edge(5054, 5055).
edge(5055, 5056).
edge(5056, 5057).
edge(5057, 5058).
edge(5058, 5059).
edge(5059, 5060).
edge(5060, 5061).
edge(5061, 5062).
edge(5062, 5063).
edge(5063, 5064).
edge(5064, 5065).
edge(5065, 5066).
edge(5066, 5067).
edge(5067, 5068).
edge(5068, 5069).
edge(5069, 5070).
edge(5070, 5071).
edge(5071, 5072).
edge(5072, 5073).
edge(5073, 5074).
edge(5074, 5075).
edge(5075, 5076).
edge(5076, 5077).
edge(5077, 5078).
edge(5078, 5079).
edge(5079, 5080).
edge(5080, 5081).
edge(5081, 5082).
edge(5082, 5083).
edge(5083, 5084).
edge(5084, 5085).
edge(5085, 5086).
edge(5086, 5087).
edge(5087, 5088).
edge(5088, 5089).
edge(5089, 5090).
edge(5090, 5091).
edge(5091, 5092).
edge(5092, 5093).
edge(5093, 5094).
edge(5094, 5095).
edge(5095, 5096).
edge(5096, 5097).
edge(5097, 5098).
edge(5098, 5099).
edge(5099, 5100).
edge(5100, 5101).
edge(5101, 5102).
edge(5102, 5103).
edge(5103, 5104).
edge(5104, 5105).
edge(5105, 5106).
edge(5106, 5107).
edge(5107, 5108).
edge(5108, 5109).
edge(5109, 5110).
edge(5110, 5111).
edge(5111, 5112).
edge(5112, 5113).
edge(5113, 5114).
edge(5114, 5115).
edge(5115, 5116).
edge(5116, 5117).
edge(5117, 5118).
edge(5118, 5119).
edge(5119, 5120).
edge(5120, 5121).
edge(5121, 5122).
edge(5122, 5123).
edge(5123, 5124).
edge(5124, 5125).
edge(5125, 5126).
edge(5126, 5127).
edge(5127, 5128).
edge(5128, 5129).
edge(5129, 5130).
edge(5130, 5131).
edge(5131, 5132).
edge(5132, 5133).
edge(5133, 5134).
edge(5134, 5135).
edge(5135, 5136).
edge(5136, 5137).
edge(5137, 5138).
edge(5138, 5139).
edge(5139, 5140).
edge(5140, 5141).
edge(5141, 5142).
edge(5142, 5143).
edge(5143, 5144).
edge(5144, 5145).
edge(5145, 5146).
edge(5146, 5147).
edge(5147, 5148).
edge(5148, 5149).
edge(5149, 5150).
edge(5150, 5151).
edge(5151, 5152).
edge(5152, 5153).
edge(5153, 5154).
edge(5154, 5155).
edge(5155, 5156).
edge(5156, 5157).
edge(5157, 5158).
edge(5158, 5159).
edge(5159, 5160).
edge(5160, 5161).
edge(5161, 5162).
edge(5162, 5163).
edge(5163, 5164).
edge(5164, 5165).
edge(5165, 5166).
edge(5166, 5167).
edge(5167, 5168).
edge(5168, 5169).
edge(5169, 5170).
edge(5170, 5171).
edge(5171, 5172).
edge(5172, 5173).
edge(5173, 5174).
edge(5174, 5175).
edge(5175, 5176).
edge(5176, 5177).
edge(5177, 5178).
edge(5178, 5179).
edge(5179, 5180).
edge(5180, 5181).
edge(5181, 5182).
edge(5182, 5183).
edge(5183, 5184).
edge(5184, 5185).
edge(5185, 5186).
edge(5186, 5187).
edge(5187, 5188).
edge(5188, 5189).
edge(5189, 5190).
edge(5190, 5191).
edge(5191, 5192).
edge(5192, 5193).
edge(5193, 5194).
edge(5194, 5195).
edge(5195, 5196).
edge(5196, 5197).
edge(5197, 5198).
edge(5198, 5199).
edge(5199, 5200).
edge(5200, 5201).
edge(5201, 5202).
edge(5202, 5203).
edge(5203, 5204).
edge(5204, 5205).
edge(5205, 5206).
edge(5206, 5207).
edge(5207, 5208).
edge(5208, 5209).
edge(5209, 5210).
edge(5210, 5211).
edge(5211, 5212).
edge(5212, 5213).
edge(5213, 5214).
edge(5214, 5215).
edge(5215, 5216).
edge(5216, 5217).
edge(5217, 5218).
edge(5218, 5219).
edge(5219, 5220).
edge(5220, 5221).
edge(5221, 5222).
edge(5222, 5223).
edge(5223, 5224).
edge(5224, 5225).
edge(5225, 5226).
edge(5226, 5227).
edge(5227, 5228).
edge(5228, 5229).
edge(5229, 5230).
edge(5230, 5231).
edge(5231, 5232).
edge(5232, 5233).
edge(5233, 5234).
edge(5234, 5235).
edge(5235, 5236).
edge(5236, 5237).
edge(5237, 5238).
edge(5238, 5239).
edge(5239, 5240).
edge(5240, 5241).
edge(5241, 5242).
edge(5242, 5243).
edge(5243, 5244).
edge(5244, 5245).
edge(5245, 5246).
edge(5246, 5247).
edge(5247, 5248).
edge(5248, 5249).
edge(5249, 5250).
edge(5250, 5251).
edge(5251, 5252).
edge(5252, 5253).
edge(5253, 5254).
edge(5254, 5255).
edge(5255, 5256).
edge(5256, 5257).
edge(5257, 5258).
edge(5258, 5259).
edge(5259, 5260).
edge(5260, 5261).
edge(5261, 5262).
edge(5262, 5263).
edge(5263, 5264).
edge(5264, 5265).
edge(5265, 5266).
edge(5266, 5267).
edge(5267, 5268).
edge(5268, 5269).
edge(5269, 5270).
edge(5270, 5271).
edge(5271, 5272).
edge(5272, 5273).
edge(5273, 5274).
edge(5274, 5275).
edge(5275, 5276).
edge(5276, 5277).
edge(5277, 5278).
edge(5278, 5279).
edge(5279, 5280).
edge(5280, 5281).
edge(5281, 5282).
edge(5282, 5283).
edge(5283, 5284).
edge(5284, 5285).
edge(5285, 5286).
edge(5286, 5287).
edge(5287, 5288).
edge(5288, 5289).
edge(5289, 5290).
edge(5290, 5291).
edge(5291, 5292).
edge(5292, 5293).
edge(5293, 5294).
edge(5294, 5295).
edge(5295, 5296).
edge(5296, 5297).
edge(5297, 5298).
edge(5298, 5299).
edge(5299, 5300).
edge(5300, 5301).
edge(5301, 5302).
edge(5302, 5303).
edge(5303, 5304).
edge(5304, 5305).
edge(5305, 5306).
edge(5306, 5307).
edge(5307, 5308).
edge(5308, 5309).
edge(5309, 5310).
edge(5310, 5311).
edge(5311, 5312).
edge(5312, 5313).
edge(5313, 5314).
edge(5314, 5315).
edge(5315, 5316).
edge(5316, 5317).
edge(5317, 5318).
edge(5318, 5319).
edge(5319, 5320).
edge(5320, 5321).
edge(5321, 5322).
edge(5322, 5323).
edge(5323, 5324).
edge(5324, 5325).
edge(5325, 5326).
edge(5326, 5327).
edge(5327, 5328).
edge(5328, 5329).
edge(5329, 5330).
edge(5330, 5331).
edge(5331, 5332).
edge(5332, 5333).
edge(5333, 5334).
edge(5334, 5335).
edge(5335, 5336).
edge(5336, 5337).
edge(5337, 5338).
edge(5338, 5339).
edge(5339, 5340).
edge(5340, 5341).
edge(5341, 5342).
edge(5342, 5343).
edge(5343, 5344).
edge(5344, 5345).
edge(5345, 5346).
edge(5346, 5347).
edge(5347, 5348).
edge(5348, 5349).
edge(5349, 5350).
edge(5350, 5351).
edge(5351, 5352).
edge(5352, 5353).
edge(5353, 5354).
edge(5354, 5355).
edge(5355, 5356).
edge(5356, 5357).
edge(5357, 5358).
edge(5358, 5359).
edge(5359, 5360).
edge(5360, 5361).
edge(5361, 5362).
edge(5362, 5363).
edge(5363, 5364).
edge(5364, 5365).
edge(5365, 5366).
edge(5366, 5367).
edge(5367, 5368).
edge(5368, 5369).
edge(5369, 5370).
edge(5370, 5371).
edge(5371, 5372).
edge(5372, 5373).
edge(5373, 5374).
edge(5374, 5375).
edge(5375, 5376).
edge(5376, 5377).
edge(5377, 5378).
edge(5378, 5379).
edge(5379, 5380).
edge(5380, 5381).
edge(5381, 5382).
edge(5382, 5383).
edge(5383, 5384).
edge(5384, 5385).
edge(5385, 5386).
edge(5386, 5387).
edge(5387, 5388).
edge(5388, 5389).
edge(5389, 5390).
edge(5390, 5391).
edge(5391, 5392).
edge(5392, 5393).
edge(5393, 5394).
edge(5394, 5395).
edge(5395, 5396).
edge(5396, 5397).
edge(5397, 5398).
edge(5398, 5399).
edge(5399, 5400).
edge(5400, 5401).
edge(5401, 5402).
edge(5402, 5403).
edge(5403, 5404).
edge(5404, 5405).
edge(5405, 5406).
edge(5406, 5407).
edge(5407, 5408).
edge(5408, 5409).
edge(5409, 5410).
edge(5410, 5411).
edge(5411, 5412).
edge(5412, 5413).
edge(5413, 5414).
edge(5414, 5415).
edge(5415, 5416).
edge(5416, 5417).
edge(5417, 5418).
edge(5418, 5419).
edge(5419, 5420).
edge(5420, 5421).
edge(5421, 5422).
edge(5422, 5423).
edge(5423, 5424).
edge(5424, 5425).
edge(5425, 5426).
edge(5426, 5427).
edge(5427, 5428).
edge(5428, 5429).
edge(5429, 5430).
edge(5430, 5431).
edge(5431, 5432).
edge(5432, 5433).
edge(5433, 5434).
edge(5434, 5435).
edge(5435, 5436).
edge(5436, 5437).
edge(5437, 5438).
edge(5438, 5439).
edge(5439, 5440).
edge(5440, 5441).
edge(5441, 5442).
edge(5442, 5443).
edge(5443, 5444).
edge(5444, 5445).
edge(5445, 5446).
edge(5446, 5447).
edge(5447, 5448).
edge(5448, 5449).
edge(5449, 5450).
edge(5450, 5451).
edge(5451, 5452).
edge(5452, 5453).
edge(5453, 5454).
edge(5454, 5455).
edge(5455, 5456).
edge(5456, 5457).
edge(5457, 5458).
edge(5458, 5459).
edge(5459, 5460).
edge(5460, 5461).
edge(5461, 5462).
edge(5462, 5463).
edge(5463, 5464).
edge(5464, 5465).
edge(5465, 5466).
edge(5466, 5467).
edge(5467, 5468).
edge(5468, 5469).
edge(5469, 5470).
edge(5470, 5471).
edge(5471, 5472).
edge(5472, 5473).
edge(5473, 5474).
edge(5474, 5475).
edge(5475, 5476).
edge(5476, 5477).
edge(5477, 5478).
edge(5478, 5479).
edge(5479, 5480).
edge(5480, 5481).
edge(5481, 5482).
edge(5482, 5483).
edge(5483, 5484).
edge(5484, 5485).
edge(5485, 5486).
edge(5486, 5487).
edge(5487, 5488).
edge(5488, 5489).
edge(5489, 5490).
edge(5490, 5491).
edge(5491, 5492).
edge(5492, 5493).
edge(5493, 5494).
edge(5494, 5495).
edge(5495, 5496).
edge(5496, 5497).
edge(5497, 5498).
edge(5498, 5499).
edge(5499, 5500).
edge(5500, 5501).
edge(5501, 5502).
edge(5502, 5503).
edge(5503, 5504).
edge(5504, 5505).
edge(5505, 5506).
edge(5506, 5507).
edge(5507, 5508).
edge(5508, 5509).
edge(5509, 5510).
edge(5510, 5511).
edge(5511, 5512).
edge(5512, 5513).
edge(5513, 5514).
edge(5514, 5515).
edge(5515, 5516).
edge(5516, 5517).
edge(5517, 5518).
edge(5518, 5519).
edge(5519, 5520).
edge(5520, 5521).
edge(5521, 5522).
edge(5522, 5523).
edge(5523, 5524).
edge(5524, 5525).
edge(5525, 5526).
edge(5526, 5527).
edge(5527, 5528).
edge(5528, 5529).
edge(5529, 5530).
edge(5530, 5531).
edge(5531, 5532).
edge(5532, 5533).
edge(5533, 5534).
edge(5534, 5535).
edge(5535, 5536).
edge(5536, 5537).
edge(5537, 5538).
edge(5538, 5539).
edge(5539, 5540).
edge(5540, 5541).
edge(5541, 5542).
edge(5542, 5543).
edge(5543, 5544).
edge(5544, 5545).
edge(5545, 5546).
edge(5546, 5547).
edge(5547, 5548).
edge(5548, 5549).
edge(5549, 5550).
edge(5550, 5551).
edge(5551, 5552).
edge(5552, 5553).
edge(5553, 5554).
edge(5554, 5555).
edge(5555, 5556).
edge(5556, 5557).
edge(5557, 5558).
edge(5558, 5559).
edge(5559, 5560).
edge(5560, 5561).
edge(5561, 5562).
edge(5562, 5563).
edge(5563, 5564).
edge(5564, 5565).
edge(5565, 5566).
edge(5566, 5567).
edge(5567, 5568).
edge(5568, 5569).
edge(5569, 5570).
edge(5570, 5571).
edge(5571, 5572).
edge(5572, 5573).
edge(5573, 5574).
edge(5574, 5575).
edge(5575, 5576).
edge(5576, 5577).
edge(5577, 5578).
edge(5578, 5579).
edge(5579, 5580).
edge(5580, 5581).
edge(5581, 5582).
edge(5582, 5583).
edge(5583, 5584).
edge(5584, 5585).
edge(5585, 5586).
edge(5586, 5587).
edge(5587, 5588).
edge(5588, 5589).
edge(5589, 5590).
edge(5590, 5591).
edge(5591, 5592).
edge(5592, 5593).
edge(5593, 5594).
edge(5594, 5595).
edge(5595, 5596).
edge(5596, 5597).
edge(5597, 5598).
edge(5598, 5599).
edge(5599, 5600).
edge(5600, 5601).
edge(5601, 5602).
edge(5602, 5603).
edge(5603, 5604).
edge(5604, 5605).
edge(5605, 5606).
edge(5606, 5607).
edge(5607, 5608).
edge(5608, 5609).
edge(5609, 5610).
edge(5610, 5611).
edge(5611, 5612).
edge(5612, 5613).
edge(5613, 5614).
edge(5614, 5615).
edge(5615, 5616).
edge(5616, 5617).
edge(5617, 5618).
edge(5618, 5619).
edge(5619, 5620).
edge(5620, 5621).
edge(5621, 5622).
edge(5622, 5623).
edge(5623, 5624).
edge(5624, 5625).
edge(5625, 5626).
edge(5626, 5627).
edge(5627, 5628).
edge(5628, 5629).
edge(5629, 5630).
edge(5630, 5631).
edge(5631, 5632).
edge(5632, 5633).
edge(5633, 5634).
edge(5634, 5635).
edge(5635, 5636).
edge(5636, 5637).
edge(5637, 5638).
edge(5638, 5639).
edge(5639, 5640).
edge(5640, 5641).
edge(5641, 5642).
edge(5642, 5643).
edge(5643, 5644).
edge(5644, 5645).
edge(5645, 5646).
edge(5646, 5647).
edge(5647, 5648).
edge(5648, 5649).
edge(5649, 5650).
edge(5650, 5651).
edge(5651, 5652).
edge(5652, 5653).
edge(5653, 5654).
edge(5654, 5655).
edge(5655, 5656).
edge(5656, 5657).
edge(5657, 5658).
edge(5658, 5659).
edge(5659, 5660).
edge(5660, 5661).
edge(5661, 5662).
edge(5662, 5663).
edge(5663, 5664).
edge(5664, 5665).
edge(5665, 5666).
edge(5666, 5667).
edge(5667, 5668).
edge(5668, 5669).
edge(5669, 5670).
edge(5670, 5671).
edge(5671, 5672).
edge(5672, 5673).
edge(5673, 5674).
edge(5674, 5675).
edge(5675, 5676).
edge(5676, 5677).
edge(5677, 5678).
edge(5678, 5679).
edge(5679, 5680).
edge(5680, 5681).
edge(5681, 5682).
edge(5682, 5683).
edge(5683, 5684).
edge(5684, 5685).
edge(5685, 5686).
edge(5686, 5687).
edge(5687, 5688).
edge(5688, 5689).
edge(5689, 5690).
edge(5690, 5691).
edge(5691, 5692).
edge(5692, 5693).
edge(5693, 5694).
edge(5694, 5695).
edge(5695, 5696).
edge(5696, 5697).
edge(5697, 5698).
edge(5698, 5699).
edge(5699, 5700).
edge(5700, 5701).
edge(5701, 5702).
edge(5702, 5703).
edge(5703, 5704).
edge(5704, 5705).
edge(5705, 5706).
edge(5706, 5707).
edge(5707, 5708).
edge(5708, 5709).
edge(5709, 5710).
edge(5710, 5711).
edge(5711, 5712).
edge(5712, 5713).
edge(5713, 5714).
edge(5714, 5715).
edge(5715, 5716).
edge(5716, 5717).
edge(5717, 5718).
edge(5718, 5719).
edge(5719, 5720).
edge(5720, 5721).
edge(5721, 5722).
edge(5722, 5723).
edge(5723, 5724).
edge(5724, 5725).
edge(5725, 5726).
edge(5726, 5727).
edge(5727, 5728).
edge(5728, 5729).
edge(5729, 5730).
edge(5730, 5731).
edge(5731, 5732).
edge(5732, 5733).
edge(5733, 5734).
edge(5734, 5735).
edge(5735, 5736).
edge(5736, 5737).
edge(5737, 5738).
edge(5738, 5739).
edge(5739, 5740).
edge(5740, 5741).
edge(5741, 5742).
edge(5742, 5743).
edge(5743, 5744).
edge(5744, 5745).
edge(5745, 5746).
edge(5746, 5747).
edge(5747, 5748).
edge(5748, 5749).
edge(5749, 5750).
edge(5750, 5751).
edge(5751, 5752).
edge(5752, 5753).
edge(5753, 5754).
edge(5754, 5755).
edge(5755, 5756).
edge(5756, 5757).
edge(5757, 5758).
edge(5758, 5759).
edge(5759, 5760).
edge(5760, 5761).
edge(5761, 5762).
edge(5762, 5763).
edge(5763, 5764).
edge(5764, 5765).
edge(5765, 5766).
edge(5766, 5767).
edge(5767, 5768).
edge(5768, 5769).
edge(5769, 5770).
edge(5770, 5771).
edge(5771, 5772).
edge(5772, 5773).
edge(5773, 5774).
edge(5774, 5775).
edge(5775, 5776).
edge(5776, 5777).
edge(5777, 5778).
edge(5778, 5779).
edge(5779, 5780).
edge(5780, 5781).
edge(5781, 5782).
edge(5782, 5783).
edge(5783, 5784).
edge(5784, 5785).
edge(5785, 5786).
edge(5786, 5787).
edge(5787, 5788).
edge(5788, 5789).
edge(5789, 5790).
edge(5790, 5791).
edge(5791, 5792).
edge(5792, 5793).
edge(5793, 5794).
edge(5794, 5795).
edge(5795, 5796).
edge(5796, 5797).
edge(5797, 5798).
edge(5798, 5799).
edge(5799, 5800).
edge(5800, 5801).
edge(5801, 5802).
edge(5802, 5803).
edge(5803, 5804).
edge(5804, 5805).
edge(5805, 5806).
edge(5806, 5807).
edge(5807, 5808).
edge(5808, 5809).
edge(5809, 5810).
edge(5810, 5811).
edge(5811, 5812).
edge(5812, 5813).
edge(5813, 5814).
edge(5814, 5815).
edge(5815, 5816).
edge(5816, 5817).
edge(5817, 5818).
edge(5818, 5819).
edge(5819, 5820).
edge(5820, 5821).
edge(5821, 5822).
edge(5822, 5823).
edge(5823, 5824).
edge(5824, 5825).
edge(5825, 5826).
edge(5826, 5827).
edge(5827, 5828).
edge(5828, 5829).
edge(5829, 5830).
edge(5830, 5831).
edge(5831, 5832).
edge(5832, 5833).
edge(5833, 5834).
edge(5834, 5835).
edge(5835, 5836).
edge(5836, 5837).
edge(5837, 5838).
edge(5838, 5839).
edge(5839, 5840).
edge(5840, 5841).
edge(5841, 5842).
edge(5842, 5843).
edge(5843, 5844).
edge(5844, 5845).
edge(5845, 5846).
edge(5846, 5847).
edge(5847, 5848).
edge(5848, 5849).
edge(5849, 5850).
edge(5850, 5851).
edge(5851, 5852).
edge(5852, 5853).
edge(5853, 5854).
edge(5854, 5855).
edge(5855, 5856).
edge(5856, 5857).
edge(5857, 5858).
edge(5858, 5859).
edge(5859, 5860).
edge(5860, 5861).
edge(5861, 5862).
edge(5862, 5863).
edge(5863, 5864).
edge(5864, 5865).
edge(5865, 5866).
edge(5866, 5867).
edge(5867, 5868).
edge(5868, 5869).
edge(5869, 5870).
edge(5870, 5871).
edge(5871, 5872).
edge(5872, 5873).
edge(5873, 5874).
edge(5874, 5875).
edge(5875, 5876).
edge(5876, 5877).
edge(5877, 5878).
edge(5878, 5879).
edge(5879, 5880).
edge(5880, 5881).
edge(5881, 5882).
edge(5882, 5883).
edge(5883, 5884).
edge(5884, 5885).
edge(5885, 5886).
edge(5886, 5887).
edge(5887, 5888).
edge(5888, 5889).
edge(5889, 5890).
edge(5890, 5891).
edge(5891, 5892).
edge(5892, 5893).
edge(5893, 5894).
edge(5894, 5895).
edge(5895, 5896).
edge(5896, 5897).
edge(5897, 5898).
edge(5898, 5899).
edge(5899, 5900).
edge(5900, 5901).
edge(5901, 5902).
edge(5902, 5903).
edge(5903, 5904).
edge(5904, 5905).
edge(5905, 5906).
edge(5906, 5907).
edge(5907, 5908).
edge(5908, 5909).
edge(5909, 5910).
edge(5910, 5911).
edge(5911, 5912).
edge(5912, 5913).
edge(5913, 5914).
edge(5914, 5915).
edge(5915, 5916).
edge(5916, 5917).
edge(5917, 5918).
edge(5918, 5919).
edge(5919, 5920).
edge(5920, 5921).
edge(5921, 5922).
edge(5922, 5923).
edge(5923, 5924).
edge(5924, 5925).
edge(5925, 5926).
edge(5926, 5927).
edge(5927, 5928).
edge(5928, 5929).
edge(5929, 5930).
edge(5930, 5931).
edge(5931, 5932).
edge(5932, 5933).
edge(5933, 5934).
edge(5934, 5935).
edge(5935, 5936).
edge(5936, 5937).
edge(5937, 5938).
edge(5938, 5939).
edge(5939, 5940).
edge(5940, 5941).
edge(5941, 5942).
edge(5942, 5943).
edge(5943, 5944).
edge(5944, 5945).
edge(5945, 5946).
edge(5946, 5947).
edge(5947, 5948).
edge(5948, 5949).
edge(5949, 5950).
edge(5950, 5951).
edge(5951, 5952).
edge(5952, 5953).
edge(5953, 5954).
edge(5954, 5955).
edge(5955, 5956).
edge(5956, 5957).
edge(5957, 5958).
edge(5958, 5959).
edge(5959, 5960).
edge(5960, 5961).
edge(5961, 5962).
edge(5962, 5963).
edge(5963, 5964).
edge(5964, 5965).
edge(5965, 5966).
edge(5966, 5967).
edge(5967, 5968).
edge(5968, 5969).
edge(5969, 5970).
edge(5970, 5971).
edge(5971, 5972).
edge(5972, 5973).
edge(5973, 5974).
edge(5974, 5975).
edge(5975, 5976).
edge(5976, 5977).
edge(5977, 5978).
edge(5978, 5979).
edge(5979, 5980).
edge(5980, 5981).
edge(5981, 5982).
edge(5982, 5983).
edge(5983, 5984).
edge(5984, 5985).
edge(5985, 5986).
edge(5986, 5987).
edge(5987, 5988).
edge(5988, 5989).
edge(5989, 5990).
edge(5990, 5991).
edge(5991, 5992).
edge(5992, 5993).
edge(5993, 5994).
edge(5994, 5995).
edge(5995, 5996).
edge(5996, 5997).
edge(5997, 5998).
edge(5998, 5999).
edge(5999, 6000).
edge(6000, 6001).
edge(6001, 6002).
edge(6002, 6003).
edge(6003, 6004).
edge(6004, 6005).
edge(6005, 6006).
edge(6006, 6007).
edge(6007, 6008).
edge(6008, 6009).
edge(6009, 6010).
edge(6010, 6011).
edge(6011, 6012).
edge(6012, 6013).
edge(6013, 6014).
edge(6014, 6015).
edge(6015, 6016).
edge(6016, 6017).
edge(6017, 6018).
edge(6018, 6019).
edge(6019, 6020).
edge(6020, 6021).
edge(6021, 6022).
edge(6022, 6023).
edge(6023, 6024).
edge(6024, 6025).
edge(6025, 6026).
edge(6026, 6027).
edge(6027, 6028).
edge(6028, 6029).
edge(6029, 6030).
edge(6030, 6031).
edge(6031, 6032).
edge(6032, 6033).
edge(6033, 6034).
edge(6034, 6035).
edge(6035, 6036).
edge(6036, 6037).
edge(6037, 6038).
edge(6038, 6039).
edge(6039, 6040).
edge(6040, 6041).
edge(6041, 6042).
edge(6042, 6043).
edge(6043, 6044).
edge(6044, 6045).
edge(6045, 6046).
edge(6046, 6047).
edge(6047, 6048).
edge(6048, 6049).
edge(6049, 6050).
edge(6050, 6051).
edge(6051, 6052).
edge(6052, 6053).
edge(6053, 6054).
edge(6054, 6055).
edge(6055, 6056).
edge(6056, 6057).
edge(6057, 6058).
edge(6058, 6059).
edge(6059, 6060).
edge(6060, 6061).
edge(6061, 6062).
edge(6062, 6063).
edge(6063, 6064).
edge(6064, 6065).
edge(6065, 6066).
edge(6066, 6067).
edge(6067, 6068).
edge(6068, 6069).
edge(6069, 6070).
edge(6070, 6071).
edge(6071, 6072).
edge(6072, 6073).
edge(6073, 6074).
edge(6074, 6075).
edge(6075, 6076).
edge(6076, 6077).
edge(6077, 6078).
edge(6078, 6079).
edge(6079, 6080).
edge(6080, 6081).
edge(6081, 6082).
edge(6082, 6083).
edge(6083, 6084).
edge(6084, 6085).
edge(6085, 6086).
edge(6086, 6087).
edge(6087, 6088).
edge(6088, 6089).
edge(6089, 6090).
edge(6090, 6091).
edge(6091, 6092).
edge(6092, 6093).
edge(6093, 6094).
edge(6094, 6095).
edge(6095, 6096).
edge(6096, 6097).
edge(6097, 6098).
edge(6098, 6099).
edge(6099, 6100).
edge(6100, 6101).
edge(6101, 6102).
edge(6102, 6103).
edge(6103, 6104).
edge(6104, 6105).
edge(6105, 6106).
edge(6106, 6107).
edge(6107, 6108).
edge(6108, 6109).
edge(6109, 6110).
edge(6110, 6111).
edge(6111, 6112).
edge(6112, 6113).
edge(6113, 6114).
edge(6114, 6115).
edge(6115, 6116).
edge(6116, 6117).
edge(6117, 6118).
edge(6118, 6119).
edge(6119, 6120).
edge(6120, 6121).
edge(6121, 6122).
edge(6122, 6123).
edge(6123, 6124).
edge(6124, 6125).
edge(6125, 6126).
edge(6126, 6127).
edge(6127, 6128).
edge(6128, 6129).
edge(6129, 6130).
edge(6130, 6131).
edge(6131, 6132).
edge(6132, 6133).
edge(6133, 6134).
edge(6134, 6135).
edge(6135, 6136).
edge(6136, 6137).
edge(6137, 6138).
edge(6138, 6139).
edge(6139, 6140).
edge(6140, 6141).
edge(6141, 6142).
edge(6142, 6143).
edge(6143, 6144).
edge(6144, 6145).
edge(6145, 6146).
edge(6146, 6147).
edge(6147, 6148).
edge(6148, 6149).
edge(6149, 6150).
edge(6150, 6151).
edge(6151, 6152).
edge(6152, 6153).
edge(6153, 6154).
edge(6154, 6155).
edge(6155, 6156).
edge(6156, 6157).
edge(6157, 6158).
edge(6158, 6159).
edge(6159, 6160).
edge(6160, 6161).
edge(6161, 6162).
edge(6162, 6163).
edge(6163, 6164).
edge(6164, 6165).
edge(6165, 6166).
edge(6166, 6167).
edge(6167, 6168).
edge(6168, 6169).
edge(6169, 6170).
edge(6170, 6171).
edge(6171, 6172).
edge(6172, 6173).
edge(6173, 6174).
edge(6174, 6175).
edge(6175, 6176).
edge(6176, 6177).
edge(6177, 6178).
edge(6178, 6179).
edge(6179, 6180).
edge(6180, 6181).
edge(6181, 6182).
edge(6182, 6183).
edge(6183, 6184).
edge(6184, 6185).
edge(6185, 6186).
edge(6186, 6187).
edge(6187, 6188).
edge(6188, 6189).
edge(6189, 6190).
edge(6190, 6191).
edge(6191, 6192).
edge(6192, 6193).
edge(6193, 6194).
edge(6194, 6195).
edge(6195, 6196).
edge(6196, 6197).
edge(6197, 6198).
edge(6198, 6199).
edge(6199, 6200).
edge(6200, 6201).
edge(6201, 6202).
edge(6202, 6203).
edge(6203, 6204).
edge(6204, 6205).
edge(6205, 6206).
edge(6206, 6207).
edge(6207, 6208).
edge(6208, 6209).
edge(6209, 6210).
edge(6210, 6211).
edge(6211, 6212).
edge(6212, 6213).
edge(6213, 6214).
edge(6214, 6215).
edge(6215, 6216).
edge(6216, 6217).
edge(6217, 6218).
edge(6218, 6219).
edge(6219, 6220).
edge(6220, 6221).
edge(6221, 6222).
edge(6222, 6223).
edge(6223, 6224).
edge(6224, 6225).
edge(6225, 6226).
edge(6226, 6227).
edge(6227, 6228).
edge(6228, 6229).
edge(6229, 6230).
edge(6230, 6231).
edge(6231, 6232).
edge(6232, 6233).
edge(6233, 6234).
edge(6234, 6235).
edge(6235, 6236).
edge(6236, 6237).
edge(6237, 6238).
edge(6238, 6239).
edge(6239, 6240).
edge(6240, 6241).
edge(6241, 6242).
edge(6242, 6243).
edge(6243, 6244).
edge(6244, 6245).
edge(6245, 6246).
edge(6246, 6247).
edge(6247, 6248).
edge(6248, 6249).
edge(6249, 6250).
edge(6250, 6251).
edge(6251, 6252).
edge(6252, 6253).
edge(6253, 6254).
edge(6254, 6255).
edge(6255, 6256).
edge(6256, 6257).
edge(6257, 6258).
edge(6258, 6259).
edge(6259, 6260).
edge(6260, 6261).
edge(6261, 6262).
edge(6262, 6263).
edge(6263, 6264).
edge(6264, 6265).
edge(6265, 6266).
edge(6266, 6267).
edge(6267, 6268).
edge(6268, 6269).
edge(6269, 6270).
edge(6270, 6271).
edge(6271, 6272).
edge(6272, 6273).
edge(6273, 6274).
edge(6274, 6275).
edge(6275, 6276).
edge(6276, 6277).
edge(6277, 6278).
edge(6278, 6279).
edge(6279, 6280).
edge(6280, 6281).
edge(6281, 6282).
edge(6282, 6283).
edge(6283, 6284).
edge(6284, 6285).
edge(6285, 6286).
edge(6286, 6287).
edge(6287, 6288).
edge(6288, 6289).
edge(6289, 6290).
edge(6290, 6291).
edge(6291, 6292).
edge(6292, 6293).
edge(6293, 6294).
edge(6294, 6295).
edge(6295, 6296).
edge(6296, 6297).
edge(6297, 6298).
edge(6298, 6299).
edge(6299, 6300).
edge(6300, 6301).
edge(6301, 6302).
edge(6302, 6303).
edge(6303, 6304).
edge(6304, 6305).
edge(6305, 6306).
edge(6306, 6307).
edge(6307, 6308).
edge(6308, 6309).
edge(6309, 6310).
edge(6310, 6311).
edge(6311, 6312).
edge(6312, 6313).
edge(6313, 6314).
edge(6314, 6315).
edge(6315, 6316).
edge(6316, 6317).
edge(6317, 6318).
edge(6318, 6319).
edge(6319, 6320).
edge(6320, 6321).
edge(6321, 6322).
edge(6322, 6323).
edge(6323, 6324).
edge(6324, 6325).
edge(6325, 6326).
edge(6326, 6327).
edge(6327, 6328).
edge(6328, 6329).
edge(6329, 6330).
edge(6330, 6331).
edge(6331, 6332).
edge(6332, 6333).
edge(6333, 6334).
edge(6334, 6335).
edge(6335, 6336).
edge(6336, 6337).
edge(6337, 6338).
edge(6338, 6339).
edge(6339, 6340).
edge(6340, 6341).
edge(6341, 6342).
edge(6342, 6343).
edge(6343, 6344).
edge(6344, 6345).
edge(6345, 6346).
edge(6346, 6347).
edge(6347, 6348).
edge(6348, 6349).
edge(6349, 6350).
edge(6350, 6351).
edge(6351, 6352).
edge(6352, 6353).
edge(6353, 6354).
edge(6354, 6355).
edge(6355, 6356).
edge(6356, 6357).
edge(6357, 6358).
edge(6358, 6359).
edge(6359, 6360).
edge(6360, 6361).
edge(6361, 6362).
edge(6362, 6363).
edge(6363, 6364).
edge(6364, 6365).
edge(6365, 6366).
edge(6366, 6367).
edge(6367, 6368).
edge(6368, 6369).
edge(6369, 6370).
edge(6370, 6371).
edge(6371, 6372).
edge(6372, 6373).
edge(6373, 6374).
edge(6374, 6375).
edge(6375, 6376).
edge(6376, 6377).
edge(6377, 6378).
edge(6378, 6379).
edge(6379, 6380).
edge(6380, 6381).
edge(6381, 6382).
edge(6382, 6383).
edge(6383, 6384).
edge(6384, 6385).
edge(6385, 6386).
edge(6386, 6387).
edge(6387, 6388).
edge(6388, 6389).
edge(6389, 6390).
edge(6390, 6391).
edge(6391, 6392).
edge(6392, 6393).
edge(6393, 6394).
edge(6394, 6395).
edge(6395, 6396).
edge(6396, 6397).
edge(6397, 6398).
edge(6398, 6399).
edge(6399, 6400).
edge(6400, 6401).
edge(6401, 6402).
edge(6402, 6403).
edge(6403, 6404).
edge(6404, 6405).
edge(6405, 6406).
edge(6406, 6407).
edge(6407, 6408).
edge(6408, 6409).
edge(6409, 6410).
edge(6410, 6411).
edge(6411, 6412).
edge(6412, 6413).
edge(6413, 6414).
edge(6414, 6415).
edge(6415, 6416).
edge(6416, 6417).
edge(6417, 6418).
edge(6418, 6419).
edge(6419, 6420).
edge(6420, 6421).
edge(6421, 6422).
edge(6422, 6423).
edge(6423, 6424).
edge(6424, 6425).
edge(6425, 6426).
edge(6426, 6427).
edge(6427, 6428).
edge(6428, 6429).
edge(6429, 6430).
edge(6430, 6431).
edge(6431, 6432).
edge(6432, 6433).
edge(6433, 6434).
edge(6434, 6435).
edge(6435, 6436).
edge(6436, 6437).
edge(6437, 6438).
edge(6438, 6439).
edge(6439, 6440).
edge(6440, 6441).
edge(6441, 6442).
edge(6442, 6443).
edge(6443, 6444).
edge(6444, 6445).
edge(6445, 6446).
edge(6446, 6447).
edge(6447, 6448).
edge(6448, 6449).
edge(6449, 6450).
edge(6450, 6451).
edge(6451, 6452).
edge(6452, 6453).
edge(6453, 6454).
edge(6454, 6455).
edge(6455, 6456).
edge(6456, 6457).
edge(6457, 6458).
edge(6458, 6459).
edge(6459, 6460).
edge(6460, 6461).
edge(6461, 6462).
edge(6462, 6463).
edge(6463, 6464).
edge(6464, 6465).
edge(6465, 6466).
edge(6466, 6467).
edge(6467, 6468).
edge(6468, 6469).
edge(6469, 6470).
edge(6470, 6471).
edge(6471, 6472).
edge(6472, 6473).
edge(6473, 6474).
edge(6474, 6475).
edge(6475, 6476).
edge(6476, 6477).
edge(6477, 6478).
edge(6478, 6479).
edge(6479, 6480).
edge(6480, 6481).
edge(6481, 6482).
edge(6482, 6483).
edge(6483, 6484).
edge(6484, 6485).
edge(6485, 6486).
edge(6486, 6487).
edge(6487, 6488).
edge(6488, 6489).
edge(6489, 6490).
edge(6490, 6491).
edge(6491, 6492).
edge(6492, 6493).
edge(6493, 6494).
edge(6494, 6495).
edge(6495, 6496).
edge(6496, 6497).
edge(6497, 6498).
edge(6498, 6499).
edge(6499, 6500).
edge(6500, 6501).
edge(6501, 6502).
edge(6502, 6503).
edge(6503, 6504).
edge(6504, 6505).
edge(6505, 6506).
edge(6506, 6507).
edge(6507, 6508).
edge(6508, 6509).
edge(6509, 6510).
edge(6510, 6511).
edge(6511, 6512).
edge(6512, 6513).
edge(6513, 6514).
edge(6514, 6515).
edge(6515, 6516).
edge(6516, 6517).
edge(6517, 6518).
edge(6518, 6519).
edge(6519, 6520).
edge(6520, 6521).
edge(6521, 6522).
edge(6522, 6523).
edge(6523, 6524).
edge(6524, 6525).
edge(6525, 6526).
edge(6526, 6527).
edge(6527, 6528).
edge(6528, 6529).
edge(6529, 6530).
edge(6530, 6531).
edge(6531, 6532).
edge(6532, 6533).
edge(6533, 6534).
edge(6534, 6535).
edge(6535, 6536).
edge(6536, 6537).
edge(6537, 6538).
edge(6538, 6539).
edge(6539, 6540).
edge(6540, 6541).
edge(6541, 6542).
edge(6542, 6543).
edge(6543, 6544).
edge(6544, 6545).
edge(6545, 6546).
edge(6546, 6547).
edge(6547, 6548).
edge(6548, 6549).
edge(6549, 6550).
edge(6550, 6551).
edge(6551, 6552).
edge(6552, 6553).
edge(6553, 6554).
edge(6554, 6555).
edge(6555, 6556).
edge(6556, 6557).
edge(6557, 6558).
edge(6558, 6559).
edge(6559, 6560).
edge(6560, 6561).
edge(6561, 6562).
edge(6562, 6563).
edge(6563, 6564).
edge(6564, 6565).
edge(6565, 6566).
edge(6566, 6567).
edge(6567, 6568).
edge(6568, 6569).
edge(6569, 6570).
edge(6570, 6571).
edge(6571, 6572).
edge(6572, 6573).
edge(6573, 6574).
edge(6574, 6575).
edge(6575, 6576).
edge(6576, 6577).
edge(6577, 6578).
edge(6578, 6579).
edge(6579, 6580).
edge(6580, 6581).
edge(6581, 6582).
edge(6582, 6583).
edge(6583, 6584).
edge(6584, 6585).
edge(6585, 6586).
edge(6586, 6587).
edge(6587, 6588).
edge(6588, 6589).
edge(6589, 6590).
edge(6590, 6591).
edge(6591, 6592).
edge(6592, 6593).
edge(6593, 6594).
edge(6594, 6595).
edge(6595, 6596).
edge(6596, 6597).
edge(6597, 6598).
edge(6598, 6599).
edge(6599, 6600).
edge(6600, 6601).
edge(6601, 6602).
edge(6602, 6603).
edge(6603, 6604).
edge(6604, 6605).
edge(6605, 6606).
edge(6606, 6607).
edge(6607, 6608).
edge(6608, 6609).
edge(6609, 6610).
edge(6610, 6611).
edge(6611, 6612).
edge(6612, 6613).
edge(6613, 6614).
edge(6614, 6615).
edge(6615, 6616).
edge(6616, 6617).
edge(6617, 6618).
edge(6618, 6619).
edge(6619, 6620).
edge(6620, 6621).
edge(6621, 6622).
edge(6622, 6623).
edge(6623, 6624).
edge(6624, 6625).
edge(6625, 6626).
edge(6626, 6627).
edge(6627, 6628).
edge(6628, 6629).
edge(6629, 6630).
edge(6630, 6631).
edge(6631, 6632).
edge(6632, 6633).
edge(6633, 6634).
edge(6634, 6635).
edge(6635, 6636).
edge(6636, 6637).
edge(6637, 6638).
edge(6638, 6639).
edge(6639, 6640).
edge(6640, 6641).
edge(6641, 6642).
edge(6642, 6643).
edge(6643, 6644).
edge(6644, 6645).
edge(6645, 6646).
edge(6646, 6647).
edge(6647, 6648).
edge(6648, 6649).
edge(6649, 6650).
edge(6650, 6651).
edge(6651, 6652).
edge(6652, 6653).
edge(6653, 6654).
edge(6654, 6655).
edge(6655, 6656).
edge(6656, 6657).
edge(6657, 6658).
edge(6658, 6659).
edge(6659, 6660).
edge(6660, 6661).
edge(6661, 6662).
edge(6662, 6663).
edge(6663, 6664).
edge(6664, 6665).
edge(6665, 6666).
edge(6666, 6667).
edge(6667, 6668).
edge(6668, 6669).
edge(6669, 6670).
edge(6670, 6671).
edge(6671, 6672).
edge(6672, 6673).
edge(6673, 6674).
edge(6674, 6675).
edge(6675, 6676).
edge(6676, 6677).
edge(6677, 6678).
edge(6678, 6679).
edge(6679, 6680).
edge(6680, 6681).
edge(6681, 6682).
edge(6682, 6683).
edge(6683, 6684).
edge(6684, 6685).
edge(6685, 6686).
edge(6686, 6687).
edge(6687, 6688).
edge(6688, 6689).
edge(6689, 6690).
edge(6690, 6691).
edge(6691, 6692).
edge(6692, 6693).
edge(6693, 6694).
edge(6694, 6695).
edge(6695, 6696).
edge(6696, 6697).
edge(6697, 6698).
edge(6698, 6699).
edge(6699, 6700).
edge(6700, 6701).
edge(6701, 6702).
edge(6702, 6703).
edge(6703, 6704).
edge(6704, 6705).
edge(6705, 6706).
edge(6706, 6707).
edge(6707, 6708).
edge(6708, 6709).
edge(6709, 6710).
edge(6710, 6711).
edge(6711, 6712).
edge(6712, 6713).
edge(6713, 6714).
edge(6714, 6715).
edge(6715, 6716).
edge(6716, 6717).
edge(6717, 6718).
edge(6718, 6719).
edge(6719, 6720).
edge(6720, 6721).
edge(6721, 6722).
edge(6722, 6723).
edge(6723, 6724).
edge(6724, 6725).
edge(6725, 6726).
edge(6726, 6727).
edge(6727, 6728).
edge(6728, 6729).
edge(6729, 6730).
edge(6730, 6731).
edge(6731, 6732).
edge(6732, 6733).
edge(6733, 6734).
edge(6734, 6735).
edge(6735, 6736).
edge(6736, 6737).
edge(6737, 6738).
edge(6738, 6739).
edge(6739, 6740).
edge(6740, 6741).
edge(6741, 6742).
edge(6742, 6743).
edge(6743, 6744).
edge(6744, 6745).
edge(6745, 6746).
edge(6746, 6747).
edge(6747, 6748).
edge(6748, 6749).
edge(6749, 6750).
edge(6750, 6751).
edge(6751, 6752).
edge(6752, 6753).
edge(6753, 6754).
edge(6754, 6755).
edge(6755, 6756).
edge(6756, 6757).
edge(6757, 6758).
edge(6758, 6759).
edge(6759, 6760).
edge(6760, 6761).
edge(6761, 6762).
edge(6762, 6763).
edge(6763, 6764).
edge(6764, 6765).
edge(6765, 6766).
edge(6766, 6767).
edge(6767, 6768).
edge(6768, 6769).
edge(6769, 6770).
edge(6770, 6771).
edge(6771, 6772).
edge(6772, 6773).
edge(6773, 6774).
edge(6774, 6775).
edge(6775, 6776).
edge(6776, 6777).
edge(6777, 6778).
edge(6778, 6779).
edge(6779, 6780).
edge(6780, 6781).
edge(6781, 6782).
edge(6782, 6783).
edge(6783, 6784).
edge(6784, 6785).
edge(6785, 6786).
edge(6786, 6787).
edge(6787, 6788).
edge(6788, 6789).
edge(6789, 6790).
edge(6790, 6791).
edge(6791, 6792).
edge(6792, 6793).
edge(6793, 6794).
edge(6794, 6795).
edge(6795, 6796).
edge(6796, 6797).
edge(6797, 6798).
edge(6798, 6799).
edge(6799, 6800).
edge(6800, 6801).
edge(6801, 6802).
edge(6802, 6803).
edge(6803, 6804).
edge(6804, 6805).
edge(6805, 6806).
edge(6806, 6807).
edge(6807, 6808).
edge(6808, 6809).
edge(6809, 6810).
edge(6810, 6811).
edge(6811, 6812).
edge(6812, 6813).
edge(6813, 6814).
edge(6814, 6815).
edge(6815, 6816).
edge(6816, 6817).
edge(6817, 6818).
edge(6818, 6819).
edge(6819, 6820).
edge(6820, 6821).
edge(6821, 6822).
edge(6822, 6823).
edge(6823, 6824).
edge(6824, 6825).
edge(6825, 6826).
edge(6826, 6827).
edge(6827, 6828).
edge(6828, 6829).
edge(6829, 6830).
edge(6830, 6831).
edge(6831, 6832).
edge(6832, 6833).
edge(6833, 6834).
edge(6834, 6835).
edge(6835, 6836).
edge(6836, 6837).
edge(6837, 6838).
edge(6838, 6839).
edge(6839, 6840).
edge(6840, 6841).
edge(6841, 6842).
edge(6842, 6843).
edge(6843, 6844).
edge(6844, 6845).
edge(6845, 6846).
edge(6846, 6847).
edge(6847, 6848).
edge(6848, 6849).
edge(6849, 6850).
edge(6850, 6851).
edge(6851, 6852).
edge(6852, 6853).
edge(6853, 6854).
edge(6854, 6855).
edge(6855, 6856).
edge(6856, 6857).
edge(6857, 6858).
edge(6858, 6859).
edge(6859, 6860).
edge(6860, 6861).
edge(6861, 6862).
edge(6862, 6863).
edge(6863, 6864).
edge(6864, 6865).
edge(6865, 6866).
edge(6866, 6867).
edge(6867, 6868).
edge(6868, 6869).
edge(6869, 6870).
edge(6870, 6871).
edge(6871, 6872).
edge(6872, 6873).
edge(6873, 6874).
edge(6874, 6875).
edge(6875, 6876).
edge(6876, 6877).
edge(6877, 6878).
edge(6878, 6879).
edge(6879, 6880).
edge(6880, 6881).
edge(6881, 6882).
edge(6882, 6883).
edge(6883, 6884).
edge(6884, 6885).
edge(6885, 6886).
edge(6886, 6887).
edge(6887, 6888).
edge(6888, 6889).
edge(6889, 6890).
edge(6890, 6891).
edge(6891, 6892).
edge(6892, 6893).
edge(6893, 6894).
edge(6894, 6895).
edge(6895, 6896).
edge(6896, 6897).
edge(6897, 6898).
edge(6898, 6899).
edge(6899, 6900).
edge(6900, 6901).
edge(6901, 6902).
edge(6902, 6903).
edge(6903, 6904).
edge(6904, 6905).
edge(6905, 6906).
edge(6906, 6907).
edge(6907, 6908).
edge(6908, 6909).
edge(6909, 6910).
edge(6910, 6911).
edge(6911, 6912).
edge(6912, 6913).
edge(6913, 6914).
edge(6914, 6915).
edge(6915, 6916).
edge(6916, 6917).
edge(6917, 6918).
edge(6918, 6919).
edge(6919, 6920).
edge(6920, 6921).
edge(6921, 6922).
edge(6922, 6923).
edge(6923, 6924).
edge(6924, 6925).
edge(6925, 6926).
edge(6926, 6927).
edge(6927, 6928).
edge(6928, 6929).
edge(6929, 6930).
edge(6930, 6931).
edge(6931, 6932).
edge(6932, 6933).
edge(6933, 6934).
edge(6934, 6935).
edge(6935, 6936).
edge(6936, 6937).
edge(6937, 6938).
edge(6938, 6939).
edge(6939, 6940).
edge(6940, 6941).
edge(6941, 6942).
edge(6942, 6943).
edge(6943, 6944).
edge(6944, 6945).
edge(6945, 6946).
edge(6946, 6947).
edge(6947, 6948).
edge(6948, 6949).
edge(6949, 6950).
edge(6950, 6951).
edge(6951, 6952).
edge(6952, 6953).
edge(6953, 6954).
edge(6954, 6955).
edge(6955, 6956).
edge(6956, 6957).
edge(6957, 6958).
edge(6958, 6959).
edge(6959, 6960).
edge(6960, 6961).
edge(6961, 6962).
edge(6962, 6963).
edge(6963, 6964).
edge(6964, 6965).
edge(6965, 6966).
edge(6966, 6967).
edge(6967, 6968).
edge(6968, 6969).
edge(6969, 6970).
edge(6970, 6971).
edge(6971, 6972).
edge(6972, 6973).
edge(6973, 6974).
edge(6974, 6975).
edge(6975, 6976).
edge(6976, 6977).
edge(6977, 6978).
edge(6978, 6979).
edge(6979, 6980).
edge(6980, 6981).
edge(6981, 6982).
edge(6982, 6983).
edge(6983, 6984).
edge(6984, 6985).
edge(6985, 6986).
edge(6986, 6987).
edge(6987, 6988).
edge(6988, 6989).
edge(6989, 6990).
edge(6990, 6991).
edge(6991, 6992).
edge(6992, 6993).
edge(6993, 6994).
edge(6994, 6995).
edge(6995, 6996).
edge(6996, 6997).
edge(6997, 6998).
edge(6998, 6999).
edge(6999, 7000).
edge(7000, 7001).
edge(7001, 7002).
edge(7002, 7003).
edge(7003, 7004).
edge(7004, 7005).
edge(7005, 7006).
edge(7006, 7007).
edge(7007, 7008).
edge(7008, 7009).
edge(7009, 7010).
edge(7010, 7011).
edge(7011, 7012).
edge(7012, 7013).
edge(7013, 7014).
edge(7014, 7015).
edge(7015, 7016).
edge(7016, 7017).
edge(7017, 7018).
edge(7018, 7019).
edge(7019, 7020).
edge(7020, 7021).
edge(7021, 7022).
edge(7022, 7023).
edge(7023, 7024).
edge(7024, 7025).
edge(7025, 7026).
edge(7026, 7027).
edge(7027, 7028).
edge(7028, 7029).
edge(7029, 7030).
edge(7030, 7031).
edge(7031, 7032).
edge(7032, 7033).
edge(7033, 7034).
edge(7034, 7035).
edge(7035, 7036).
edge(7036, 7037).
edge(7037, 7038).
edge(7038, 7039).
edge(7039, 7040).
edge(7040, 7041).
edge(7041, 7042).
edge(7042, 7043).
edge(7043, 7044).
edge(7044, 7045).
edge(7045, 7046).
edge(7046, 7047).
edge(7047, 7048).
edge(7048, 7049).
edge(7049, 7050).
edge(7050, 7051).
edge(7051, 7052).
edge(7052, 7053).
edge(7053, 7054).
edge(7054, 7055).
edge(7055, 7056).
edge(7056, 7057).
edge(7057, 7058).
edge(7058, 7059).
edge(7059, 7060).
edge(7060, 7061).
edge(7061, 7062).
edge(7062, 7063).
edge(7063, 7064).
edge(7064, 7065).
edge(7065, 7066).
edge(7066, 7067).
edge(7067, 7068).
edge(7068, 7069).
edge(7069, 7070).
edge(7070, 7071).
edge(7071, 7072).
edge(7072, 7073).
edge(7073, 7074).
edge(7074, 7075).
edge(7075, 7076).
edge(7076, 7077).
edge(7077, 7078).
edge(7078, 7079).
edge(7079, 7080).
edge(7080, 7081).
edge(7081, 7082).
edge(7082, 7083).
edge(7083, 7084).
edge(7084, 7085).
edge(7085, 7086).
edge(7086, 7087).
edge(7087, 7088).
edge(7088, 7089).
edge(7089, 7090).
edge(7090, 7091).
edge(7091, 7092).
edge(7092, 7093).
edge(7093, 7094).
edge(7094, 7095).
edge(7095, 7096).
edge(7096, 7097).
edge(7097, 7098).
edge(7098, 7099).
edge(7099, 7100).
edge(7100, 7101).
edge(7101, 7102).
edge(7102, 7103).
edge(7103, 7104).
edge(7104, 7105).
edge(7105, 7106).
edge(7106, 7107).
edge(7107, 7108).
edge(7108, 7109).
edge(7109, 7110).
edge(7110, 7111).
edge(7111, 7112).
edge(7112, 7113).
edge(7113, 7114).
edge(7114, 7115).
edge(7115, 7116).
edge(7116, 7117).
edge(7117, 7118).
edge(7118, 7119).
edge(7119, 7120).
edge(7120, 7121).
edge(7121, 7122).
edge(7122, 7123).
edge(7123, 7124).
edge(7124, 7125).
edge(7125, 7126).
edge(7126, 7127).
edge(7127, 7128).
edge(7128, 7129).
edge(7129, 7130).
edge(7130, 7131).
edge(7131, 7132).
edge(7132, 7133).
edge(7133, 7134).
edge(7134, 7135).
edge(7135, 7136).
edge(7136, 7137).
edge(7137, 7138).
edge(7138, 7139).
edge(7139, 7140).
edge(7140, 7141).
edge(7141, 7142).
edge(7142, 7143).
edge(7143, 7144).
edge(7144, 7145).
edge(7145, 7146).
edge(7146, 7147).
edge(7147, 7148).
edge(7148, 7149).
edge(7149, 7150).
edge(7150, 7151).
edge(7151, 7152).
edge(7152, 7153).
edge(7153, 7154).
edge(7154, 7155).
edge(7155, 7156).
edge(7156, 7157).
edge(7157, 7158).
edge(7158, 7159).
edge(7159, 7160).
edge(7160, 7161).
edge(7161, 7162).
edge(7162, 7163).
edge(7163, 7164).
edge(7164, 7165).
edge(7165, 7166).
edge(7166, 7167).
edge(7167, 7168).
edge(7168, 7169).
edge(7169, 7170).
edge(7170, 7171).
edge(7171, 7172).
edge(7172, 7173).
edge(7173, 7174).
edge(7174, 7175).
edge(7175, 7176).
edge(7176, 7177).
edge(7177, 7178).
edge(7178, 7179).
edge(7179, 7180).
edge(7180, 7181).
edge(7181, 7182).
edge(7182, 7183).
edge(7183, 7184).
edge(7184, 7185).
edge(7185, 7186).
edge(7186, 7187).
edge(7187, 7188).
edge(7188, 7189).
edge(7189, 7190).
edge(7190, 7191).
edge(7191, 7192).
edge(7192, 7193).
edge(7193, 7194).
edge(7194, 7195).
edge(7195, 7196).
edge(7196, 7197).
edge(7197, 7198).
edge(7198, 7199).
edge(7199, 7200).
edge(7200, 7201).
edge(7201, 7202).
edge(7202, 7203).
edge(7203, 7204).
edge(7204, 7205).
edge(7205, 7206).
edge(7206, 7207).
edge(7207, 7208).
edge(7208, 7209).
edge(7209, 7210).
edge(7210, 7211).
edge(7211, 7212).
edge(7212, 7213).
edge(7213, 7214).
edge(7214, 7215).
edge(7215, 7216).
edge(7216, 7217).
edge(7217, 7218).
edge(7218, 7219).
edge(7219, 7220).
edge(7220, 7221).
edge(7221, 7222).
edge(7222, 7223).
edge(7223, 7224).
edge(7224, 7225).
edge(7225, 7226).
edge(7226, 7227).
edge(7227, 7228).
edge(7228, 7229).
edge(7229, 7230).
edge(7230, 7231).
edge(7231, 7232).
edge(7232, 7233).
edge(7233, 7234).
edge(7234, 7235).
edge(7235, 7236).
edge(7236, 7237).
edge(7237, 7238).
edge(7238, 7239).
edge(7239, 7240).
edge(7240, 7241).
edge(7241, 7242).
edge(7242, 7243).
edge(7243, 7244).
edge(7244, 7245).
edge(7245, 7246).
edge(7246, 7247).
edge(7247, 7248).
edge(7248, 7249).
edge(7249, 7250).
edge(7250, 7251).
edge(7251, 7252).
edge(7252, 7253).
edge(7253, 7254).
edge(7254, 7255).
edge(7255, 7256).
edge(7256, 7257).
edge(7257, 7258).
edge(7258, 7259).
edge(7259, 7260).
edge(7260, 7261).
edge(7261, 7262).
edge(7262, 7263).
edge(7263, 7264).
edge(7264, 7265).
edge(7265, 7266).
edge(7266, 7267).
edge(7267, 7268).
edge(7268, 7269).
edge(7269, 7270).
edge(7270, 7271).
edge(7271, 7272).
edge(7272, 7273).
edge(7273, 7274).
edge(7274, 7275).
edge(7275, 7276).
edge(7276, 7277).
edge(7277, 7278).
edge(7278, 7279).
edge(7279, 7280).
edge(7280, 7281).
edge(7281, 7282).
edge(7282, 7283).
edge(7283, 7284).
edge(7284, 7285).
edge(7285, 7286).
edge(7286, 7287).
edge(7287, 7288).
edge(7288, 7289).
edge(7289, 7290).
edge(7290, 7291).
edge(7291, 7292).
edge(7292, 7293).
edge(7293, 7294).
edge(7294, 7295).
edge(7295, 7296).
edge(7296, 7297).
edge(7297, 7298).
edge(7298, 7299).
edge(7299, 7300).
edge(7300, 7301).
edge(7301, 7302).
edge(7302, 7303).
edge(7303, 7304).
edge(7304, 7305).
edge(7305, 7306).
edge(7306, 7307).
edge(7307, 7308).
edge(7308, 7309).
edge(7309, 7310).
edge(7310, 7311).
edge(7311, 7312).
edge(7312, 7313).
edge(7313, 7314).
edge(7314, 7315).
edge(7315, 7316).
edge(7316, 7317).
edge(7317, 7318).
edge(7318, 7319).
edge(7319, 7320).
edge(7320, 7321).
edge(7321, 7322).
edge(7322, 7323).
edge(7323, 7324).
edge(7324, 7325).
edge(7325, 7326).
edge(7326, 7327).
edge(7327, 7328).
edge(7328, 7329).
edge(7329, 7330).
edge(7330, 7331).
edge(7331, 7332).
edge(7332, 7333).
edge(7333, 7334).
edge(7334, 7335).
edge(7335, 7336).
edge(7336, 7337).
edge(7337, 7338).
edge(7338, 7339).
edge(7339, 7340).
edge(7340, 7341).
edge(7341, 7342).
edge(7342, 7343).
edge(7343, 7344).
edge(7344, 7345).
edge(7345, 7346).
edge(7346, 7347).
edge(7347, 7348).
edge(7348, 7349).
edge(7349, 7350).
edge(7350, 7351).
edge(7351, 7352).
edge(7352, 7353).
edge(7353, 7354).
edge(7354, 7355).
edge(7355, 7356).
edge(7356, 7357).
edge(7357, 7358).
edge(7358, 7359).
edge(7359, 7360).
edge(7360, 7361).
edge(7361, 7362).
edge(7362, 7363).
edge(7363, 7364).
edge(7364, 7365).
edge(7365, 7366).
edge(7366, 7367).
edge(7367, 7368).
edge(7368, 7369).
edge(7369, 7370).
edge(7370, 7371).
edge(7371, 7372).
edge(7372, 7373).
edge(7373, 7374).
edge(7374, 7375).
edge(7375, 7376).
edge(7376, 7377).
edge(7377, 7378).
edge(7378, 7379).
edge(7379, 7380).
edge(7380, 7381).
edge(7381, 7382).
edge(7382, 7383).
edge(7383, 7384).
edge(7384, 7385).
edge(7385, 7386).
edge(7386, 7387).
edge(7387, 7388).
edge(7388, 7389).
edge(7389, 7390).
edge(7390, 7391).
edge(7391, 7392).
edge(7392, 7393).
edge(7393, 7394).
edge(7394, 7395).
edge(7395, 7396).
edge(7396, 7397).
edge(7397, 7398).
edge(7398, 7399).
edge(7399, 7400).
edge(7400, 7401).
edge(7401, 7402).
edge(7402, 7403).
edge(7403, 7404).
edge(7404, 7405).
edge(7405, 7406).
edge(7406, 7407).
edge(7407, 7408).
edge(7408, 7409).
edge(7409, 7410).
edge(7410, 7411).
edge(7411, 7412).
edge(7412, 7413).
edge(7413, 7414).
edge(7414, 7415).
edge(7415, 7416).
edge(7416, 7417).
edge(7417, 7418).
edge(7418, 7419).
edge(7419, 7420).
edge(7420, 7421).
edge(7421, 7422).
edge(7422, 7423).
edge(7423, 7424).
edge(7424, 7425).
edge(7425, 7426).
edge(7426, 7427).
edge(7427, 7428).
edge(7428, 7429).
edge(7429, 7430).
edge(7430, 7431).
edge(7431, 7432).
edge(7432, 7433).
edge(7433, 7434).
edge(7434, 7435).
edge(7435, 7436).
edge(7436, 7437).
edge(7437, 7438).
edge(7438, 7439).
edge(7439, 7440).
edge(7440, 7441).
edge(7441, 7442).
edge(7442, 7443).
edge(7443, 7444).
edge(7444, 7445).
edge(7445, 7446).
edge(7446, 7447).
edge(7447, 7448).
edge(7448, 7449).
edge(7449, 7450).
edge(7450, 7451).
edge(7451, 7452).
edge(7452, 7453).
edge(7453, 7454).
edge(7454, 7455).
edge(7455, 7456).
edge(7456, 7457).
edge(7457, 7458).
edge(7458, 7459).
edge(7459, 7460).
edge(7460, 7461).
edge(7461, 7462).
edge(7462, 7463).
edge(7463, 7464).
edge(7464, 7465).
edge(7465, 7466).
edge(7466, 7467).
edge(7467, 7468).
edge(7468, 7469).
edge(7469, 7470).
edge(7470, 7471).
edge(7471, 7472).
edge(7472, 7473).
edge(7473, 7474).
edge(7474, 7475).
edge(7475, 7476).
edge(7476, 7477).
edge(7477, 7478).
edge(7478, 7479).
edge(7479, 7480).
edge(7480, 7481).
edge(7481, 7482).
edge(7482, 7483).
edge(7483, 7484).
edge(7484, 7485).
edge(7485, 7486).
edge(7486, 7487).
edge(7487, 7488).
edge(7488, 7489).
edge(7489, 7490).
edge(7490, 7491).
edge(7491, 7492).
edge(7492, 7493).
edge(7493, 7494).
edge(7494, 7495).
edge(7495, 7496).
edge(7496, 7497).
edge(7497, 7498).
edge(7498, 7499).
edge(7499, 7500).
edge(7500, 7501).
edge(7501, 7502).
edge(7502, 7503).
edge(7503, 7504).
edge(7504, 7505).
edge(7505, 7506).
edge(7506, 7507).
edge(7507, 7508).
edge(7508, 7509).
edge(7509, 7510).
edge(7510, 7511).
edge(7511, 7512).
edge(7512, 7513).
edge(7513, 7514).
edge(7514, 7515).
edge(7515, 7516).
edge(7516, 7517).
edge(7517, 7518).
edge(7518, 7519).
edge(7519, 7520).
edge(7520, 7521).
edge(7521, 7522).
edge(7522, 7523).
edge(7523, 7524).
edge(7524, 7525).
edge(7525, 7526).
edge(7526, 7527).
edge(7527, 7528).
edge(7528, 7529).
edge(7529, 7530).
edge(7530, 7531).
edge(7531, 7532).
edge(7532, 7533).
edge(7533, 7534).
edge(7534, 7535).
edge(7535, 7536).
edge(7536, 7537).
edge(7537, 7538).
edge(7538, 7539).
edge(7539, 7540).
edge(7540, 7541).
edge(7541, 7542).
edge(7542, 7543).
edge(7543, 7544).
edge(7544, 7545).
edge(7545, 7546).
edge(7546, 7547).
edge(7547, 7548).
edge(7548, 7549).
edge(7549, 7550).
edge(7550, 7551).
edge(7551, 7552).
edge(7552, 7553).
edge(7553, 7554).
edge(7554, 7555).
edge(7555, 7556).
edge(7556, 7557).
edge(7557, 7558).
edge(7558, 7559).
edge(7559, 7560).
edge(7560, 7561).
edge(7561, 7562).
edge(7562, 7563).
edge(7563, 7564).
edge(7564, 7565).
edge(7565, 7566).
edge(7566, 7567).
edge(7567, 7568).
edge(7568, 7569).
edge(7569, 7570).
edge(7570, 7571).
edge(7571, 7572).
edge(7572, 7573).
edge(7573, 7574).
edge(7574, 7575).
edge(7575, 7576).
edge(7576, 7577).
edge(7577, 7578).
edge(7578, 7579).
edge(7579, 7580).
edge(7580, 7581).
edge(7581, 7582).
edge(7582, 7583).
edge(7583, 7584).
edge(7584, 7585).
edge(7585, 7586).
edge(7586, 7587).
edge(7587, 7588).
edge(7588, 7589).
edge(7589, 7590).
edge(7590, 7591).
edge(7591, 7592).
edge(7592, 7593).
edge(7593, 7594).
edge(7594, 7595).
edge(7595, 7596).
edge(7596, 7597).
edge(7597, 7598).
edge(7598, 7599).
edge(7599, 7600).
edge(7600, 7601).
edge(7601, 7602).
edge(7602, 7603).
edge(7603, 7604).
edge(7604, 7605).
edge(7605, 7606).
edge(7606, 7607).
edge(7607, 7608).
edge(7608, 7609).
edge(7609, 7610).
edge(7610, 7611).
edge(7611, 7612).
edge(7612, 7613).
edge(7613, 7614).
edge(7614, 7615).
edge(7615, 7616).
edge(7616, 7617).
edge(7617, 7618).
edge(7618, 7619).
edge(7619, 7620).
edge(7620, 7621).
edge(7621, 7622).
edge(7622, 7623).
edge(7623, 7624).
edge(7624, 7625).
edge(7625, 7626).
edge(7626, 7627).
edge(7627, 7628).
edge(7628, 7629).
edge(7629, 7630).
edge(7630, 7631).
edge(7631, 7632).
edge(7632, 7633).
edge(7633, 7634).
edge(7634, 7635).
edge(7635, 7636).
edge(7636, 7637).
edge(7637, 7638).
edge(7638, 7639).
edge(7639, 7640).
edge(7640, 7641).
edge(7641, 7642).
edge(7642, 7643).
edge(7643, 7644).
edge(7644, 7645).
edge(7645, 7646).
edge(7646, 7647).
edge(7647, 7648).
edge(7648, 7649).
edge(7649, 7650).
edge(7650, 7651).
edge(7651, 7652).
edge(7652, 7653).
edge(7653, 7654).
edge(7654, 7655).
edge(7655, 7656).
edge(7656, 7657).
edge(7657, 7658).
edge(7658, 7659).
edge(7659, 7660).
edge(7660, 7661).
edge(7661, 7662).
edge(7662, 7663).
edge(7663, 7664).
edge(7664, 7665).
edge(7665, 7666).
edge(7666, 7667).
edge(7667, 7668).
edge(7668, 7669).
edge(7669, 7670).
edge(7670, 7671).
edge(7671, 7672).
edge(7672, 7673).
edge(7673, 7674).
edge(7674, 7675).
edge(7675, 7676).
edge(7676, 7677).
edge(7677, 7678).
edge(7678, 7679).
edge(7679, 7680).
edge(7680, 7681).
edge(7681, 7682).
edge(7682, 7683).
edge(7683, 7684).
edge(7684, 7685).
edge(7685, 7686).
edge(7686, 7687).
edge(7687, 7688).
edge(7688, 7689).
edge(7689, 7690).
edge(7690, 7691).
edge(7691, 7692).
edge(7692, 7693).
edge(7693, 7694).
edge(7694, 7695).
edge(7695, 7696).
edge(7696, 7697).
edge(7697, 7698).
edge(7698, 7699).
edge(7699, 7700).
edge(7700, 7701).
edge(7701, 7702).
edge(7702, 7703).
edge(7703, 7704).
edge(7704, 7705).
edge(7705, 7706).
edge(7706, 7707).
edge(7707, 7708).
edge(7708, 7709).
edge(7709, 7710).
edge(7710, 7711).
edge(7711, 7712).
edge(7712, 7713).
edge(7713, 7714).
edge(7714, 7715).
edge(7715, 7716).
edge(7716, 7717).
edge(7717, 7718).
edge(7718, 7719).
edge(7719, 7720).
edge(7720, 7721).
edge(7721, 7722).
edge(7722, 7723).
edge(7723, 7724).
edge(7724, 7725).
edge(7725, 7726).
edge(7726, 7727).
edge(7727, 7728).
edge(7728, 7729).
edge(7729, 7730).
edge(7730, 7731).
edge(7731, 7732).
edge(7732, 7733).
edge(7733, 7734).
edge(7734, 7735).
edge(7735, 7736).
edge(7736, 7737).
edge(7737, 7738).
edge(7738, 7739).
edge(7739, 7740).
edge(7740, 7741).
edge(7741, 7742).
edge(7742, 7743).
edge(7743, 7744).
edge(7744, 7745).
edge(7745, 7746).
edge(7746, 7747).
edge(7747, 7748).
edge(7748, 7749).
edge(7749, 7750).
edge(7750, 7751).
edge(7751, 7752).
edge(7752, 7753).
edge(7753, 7754).
edge(7754, 7755).
edge(7755, 7756).
edge(7756, 7757).
edge(7757, 7758).
edge(7758, 7759).
edge(7759, 7760).
edge(7760, 7761).
edge(7761, 7762).
edge(7762, 7763).
edge(7763, 7764).
edge(7764, 7765).
edge(7765, 7766).
edge(7766, 7767).
edge(7767, 7768).
edge(7768, 7769).
edge(7769, 7770).
edge(7770, 7771).
edge(7771, 7772).
edge(7772, 7773).
edge(7773, 7774).
edge(7774, 7775).
edge(7775, 7776).
edge(7776, 7777).
edge(7777, 7778).
edge(7778, 7779).
edge(7779, 7780).
edge(7780, 7781).
edge(7781, 7782).
edge(7782, 7783).
edge(7783, 7784).
edge(7784, 7785).
edge(7785, 7786).
edge(7786, 7787).
edge(7787, 7788).
edge(7788, 7789).
edge(7789, 7790).
edge(7790, 7791).
edge(7791, 7792).
edge(7792, 7793).
edge(7793, 7794).
edge(7794, 7795).
edge(7795, 7796).
edge(7796, 7797).
edge(7797, 7798).
edge(7798, 7799).
edge(7799, 7800).
edge(7800, 7801).
edge(7801, 7802).
edge(7802, 7803).
edge(7803, 7804).
edge(7804, 7805).
edge(7805, 7806).
edge(7806, 7807).
edge(7807, 7808).
edge(7808, 7809).
edge(7809, 7810).
edge(7810, 7811).
edge(7811, 7812).
edge(7812, 7813).
edge(7813, 7814).
edge(7814, 7815).
edge(7815, 7816).
edge(7816, 7817).
edge(7817, 7818).
edge(7818, 7819).
edge(7819, 7820).
edge(7820, 7821).
edge(7821, 7822).
edge(7822, 7823).
edge(7823, 7824).
edge(7824, 7825).
edge(7825, 7826).
edge(7826, 7827).
edge(7827, 7828).
edge(7828, 7829).
edge(7829, 7830).
edge(7830, 7831).
edge(7831, 7832).
edge(7832, 7833).
edge(7833, 7834).
edge(7834, 7835).
edge(7835, 7836).
edge(7836, 7837).
edge(7837, 7838).
edge(7838, 7839).
edge(7839, 7840).
edge(7840, 7841).
edge(7841, 7842).
edge(7842, 7843).
edge(7843, 7844).
edge(7844, 7845).
edge(7845, 7846).
edge(7846, 7847).
edge(7847, 7848).
edge(7848, 7849).
edge(7849, 7850).
edge(7850, 7851).
edge(7851, 7852).
edge(7852, 7853).
edge(7853, 7854).
edge(7854, 7855).
edge(7855, 7856).
edge(7856, 7857).
edge(7857, 7858).
edge(7858, 7859).
edge(7859, 7860).
edge(7860, 7861).
edge(7861, 7862).
edge(7862, 7863).
edge(7863, 7864).
edge(7864, 7865).
edge(7865, 7866).
edge(7866, 7867).
edge(7867, 7868).
edge(7868, 7869).
edge(7869, 7870).
edge(7870, 7871).
edge(7871, 7872).
edge(7872, 7873).
edge(7873, 7874).
edge(7874, 7875).
edge(7875, 7876).
edge(7876, 7877).
edge(7877, 7878).
edge(7878, 7879).
edge(7879, 7880).
edge(7880, 7881).
edge(7881, 7882).
edge(7882, 7883).
edge(7883, 7884).
edge(7884, 7885).
edge(7885, 7886).
edge(7886, 7887).
edge(7887, 7888).
edge(7888, 7889).
edge(7889, 7890).
edge(7890, 7891).
edge(7891, 7892).
edge(7892, 7893).
edge(7893, 7894).
edge(7894, 7895).
edge(7895, 7896).
edge(7896, 7897).
edge(7897, 7898).
edge(7898, 7899).
edge(7899, 7900).
edge(7900, 7901).
edge(7901, 7902).
edge(7902, 7903).
edge(7903, 7904).
edge(7904, 7905).
edge(7905, 7906).
edge(7906, 7907).
edge(7907, 7908).
edge(7908, 7909).
edge(7909, 7910).
edge(7910, 7911).
edge(7911, 7912).
edge(7912, 7913).
edge(7913, 7914).
edge(7914, 7915).
edge(7915, 7916).
edge(7916, 7917).
edge(7917, 7918).
edge(7918, 7919).
edge(7919, 7920).
edge(7920, 7921).
edge(7921, 7922).
edge(7922, 7923).
edge(7923, 7924).
edge(7924, 7925).
edge(7925, 7926).
edge(7926, 7927).
edge(7927, 7928).
edge(7928, 7929).
edge(7929, 7930).
edge(7930, 7931).
edge(7931, 7932).
edge(7932, 7933).
edge(7933, 7934).
edge(7934, 7935).
edge(7935, 7936).
edge(7936, 7937).
edge(7937, 7938).
edge(7938, 7939).
edge(7939, 7940).
edge(7940, 7941).
edge(7941, 7942).
edge(7942, 7943).
edge(7943, 7944).
edge(7944, 7945).
edge(7945, 7946).
edge(7946, 7947).
edge(7947, 7948).
edge(7948, 7949).
edge(7949, 7950).
edge(7950, 7951).
edge(7951, 7952).
edge(7952, 7953).
edge(7953, 7954).
edge(7954, 7955).
edge(7955, 7956).
edge(7956, 7957).
edge(7957, 7958).
edge(7958, 7959).
edge(7959, 7960).
edge(7960, 7961).
edge(7961, 7962).
edge(7962, 7963).
edge(7963, 7964).
edge(7964, 7965).
edge(7965, 7966).
edge(7966, 7967).
edge(7967, 7968).
edge(7968, 7969).
edge(7969, 7970).
edge(7970, 7971).
edge(7971, 7972).
edge(7972, 7973).
edge(7973, 7974).
edge(7974, 7975).
edge(7975, 7976).
edge(7976, 7977).
edge(7977, 7978).
edge(7978, 7979).
edge(7979, 7980).
edge(7980, 7981).
edge(7981, 7982).
edge(7982, 7983).
edge(7983, 7984).
edge(7984, 7985).
edge(7985, 7986).
edge(7986, 7987).
edge(7987, 7988).
edge(7988, 7989).
edge(7989, 7990).
edge(7990, 7991).
edge(7991, 7992).
edge(7992, 7993).
edge(7993, 7994).
edge(7994, 7995).
edge(7995, 7996).
edge(7996, 7997).
edge(7997, 7998).
edge(7998, 7999).
edge(7999, 8000).
edge(8000, 8001).
edge(8001, 8002).
edge(8002, 8003).
edge(8003, 8004).
edge(8004, 8005).
edge(8005, 8006).
edge(8006, 8007).
edge(8007, 8008).
edge(8008, 8009).
edge(8009, 8010).
edge(8010, 8011).
edge(8011, 8012).
edge(8012, 8013).
edge(8013, 8014).
edge(8014, 8015).
edge(8015, 8016).
edge(8016, 8017).
edge(8017, 8018).
edge(8018, 8019).
edge(8019, 8020).
edge(8020, 8021).
edge(8021, 8022).
edge(8022, 8023).
edge(8023, 8024).
edge(8024, 8025).
edge(8025, 8026).
edge(8026, 8027).
edge(8027, 8028).
edge(8028, 8029).
edge(8029, 8030).
edge(8030, 8031).
edge(8031, 8032).
edge(8032, 8033).
edge(8033, 8034).
edge(8034, 8035).
edge(8035, 8036).
edge(8036, 8037).
edge(8037, 8038).
edge(8038, 8039).
edge(8039, 8040).
edge(8040, 8041).
edge(8041, 8042).
edge(8042, 8043).
edge(8043, 8044).
edge(8044, 8045).
edge(8045, 8046).
edge(8046, 8047).
edge(8047, 8048).
edge(8048, 8049).
edge(8049, 8050).
edge(8050, 8051).
edge(8051, 8052).
edge(8052, 8053).
edge(8053, 8054).
edge(8054, 8055).
edge(8055, 8056).
edge(8056, 8057).
edge(8057, 8058).
edge(8058, 8059).
edge(8059, 8060).
edge(8060, 8061).
edge(8061, 8062).
edge(8062, 8063).
edge(8063, 8064).
edge(8064, 8065).
edge(8065, 8066).
edge(8066, 8067).
edge(8067, 8068).
edge(8068, 8069).
edge(8069, 8070).
edge(8070, 8071).
edge(8071, 8072).
edge(8072, 8073).
edge(8073, 8074).
edge(8074, 8075).
edge(8075, 8076).
edge(8076, 8077).
edge(8077, 8078).
edge(8078, 8079).
edge(8079, 8080).
edge(8080, 8081).
edge(8081, 8082).
edge(8082, 8083).
edge(8083, 8084).
edge(8084, 8085).
edge(8085, 8086).
edge(8086, 8087).
edge(8087, 8088).
edge(8088, 8089).
edge(8089, 8090).
edge(8090, 8091).
edge(8091, 8092).
edge(8092, 8093).
edge(8093, 8094).
edge(8094, 8095).
edge(8095, 8096).
edge(8096, 8097).
edge(8097, 8098).
edge(8098, 8099).
edge(8099, 8100).
edge(8100, 8101).
edge(8101, 8102).
edge(8102, 8103).
edge(8103, 8104).
edge(8104, 8105).
edge(8105, 8106).
edge(8106, 8107).
edge(8107, 8108).
edge(8108, 8109).
edge(8109, 8110).
edge(8110, 8111).
edge(8111, 8112).
edge(8112, 8113).
edge(8113, 8114).
edge(8114, 8115).
edge(8115, 8116).
edge(8116, 8117).
edge(8117, 8118).
edge(8118, 8119).
edge(8119, 8120).
edge(8120, 8121).
edge(8121, 8122).
edge(8122, 8123).
edge(8123, 8124).
edge(8124, 8125).
edge(8125, 8126).
edge(8126, 8127).
edge(8127, 8128).
edge(8128, 8129).
edge(8129, 8130).
edge(8130, 8131).
edge(8131, 8132).
edge(8132, 8133).
edge(8133, 8134).
edge(8134, 8135).
edge(8135, 8136).
edge(8136, 8137).
edge(8137, 8138).
edge(8138, 8139).
edge(8139, 8140).
edge(8140, 8141).
edge(8141, 8142).
edge(8142, 8143).
edge(8143, 8144).
edge(8144, 8145).
edge(8145, 8146).
edge(8146, 8147).
edge(8147, 8148).
edge(8148, 8149).
edge(8149, 8150).
edge(8150, 8151).
edge(8151, 8152).
edge(8152, 8153).
edge(8153, 8154).
edge(8154, 8155).
edge(8155, 8156).
edge(8156, 8157).
edge(8157, 8158).
edge(8158, 8159).
edge(8159, 8160).
edge(8160, 8161).
edge(8161, 8162).
edge(8162, 8163).
edge(8163, 8164).
edge(8164, 8165).
edge(8165, 8166).
edge(8166, 8167).
edge(8167, 8168).
edge(8168, 8169).
edge(8169, 8170).
edge(8170, 8171).
edge(8171, 8172).
edge(8172, 8173).
edge(8173, 8174).
edge(8174, 8175).
edge(8175, 8176).
edge(8176, 8177).
edge(8177, 8178).
edge(8178, 8179).
edge(8179, 8180).
edge(8180, 8181).
edge(8181, 8182).
edge(8182, 8183).
edge(8183, 8184).
edge(8184, 8185).
edge(8185, 8186).
edge(8186, 8187).
edge(8187, 8188).
edge(8188, 8189).
edge(8189, 8190).
edge(8190, 8191).
edge(8191, 8192).
edge(8192, 8193).
edge(8193, 8194).
edge(8194, 8195).
edge(8195, 8196).
edge(8196, 8197).
edge(8197, 8198).
edge(8198, 8199).
edge(8199, 8200).
edge(8200, 8201).
edge(8201, 8202).
edge(8202, 8203).
edge(8203, 8204).
edge(8204, 8205).
edge(8205, 8206).
edge(8206, 8207).
edge(8207, 8208).
edge(8208, 8209).
edge(8209, 8210).
edge(8210, 8211).
edge(8211, 8212).
edge(8212, 8213).
edge(8213, 8214).
edge(8214, 8215).
edge(8215, 8216).
edge(8216, 8217).
edge(8217, 8218).
edge(8218, 8219).
edge(8219, 8220).
edge(8220, 8221).
edge(8221, 8222).
edge(8222, 8223).
edge(8223, 8224).
edge(8224, 8225).
edge(8225, 8226).
edge(8226, 8227).
edge(8227, 8228).
edge(8228, 8229).
edge(8229, 8230).
edge(8230, 8231).
edge(8231, 8232).
edge(8232, 8233).
edge(8233, 8234).
edge(8234, 8235).
edge(8235, 8236).
edge(8236, 8237).
edge(8237, 8238).
edge(8238, 8239).
edge(8239, 8240).
edge(8240, 8241).
edge(8241, 8242).
edge(8242, 8243).
edge(8243, 8244).
edge(8244, 8245).
edge(8245, 8246).
edge(8246, 8247).
edge(8247, 8248).
edge(8248, 8249).
edge(8249, 8250).
edge(8250, 8251).
edge(8251, 8252).
edge(8252, 8253).
edge(8253, 8254).
edge(8254, 8255).
edge(8255, 8256).
edge(8256, 8257).
edge(8257, 8258).
edge(8258, 8259).
edge(8259, 8260).
edge(8260, 8261).
edge(8261, 8262).
edge(8262, 8263).
edge(8263, 8264).
edge(8264, 8265).
edge(8265, 8266).
edge(8266, 8267).
edge(8267, 8268).
edge(8268, 8269).
edge(8269, 8270).
edge(8270, 8271).
edge(8271, 8272).
edge(8272, 8273).
edge(8273, 8274).
edge(8274, 8275).
edge(8275, 8276).
edge(8276, 8277).
edge(8277, 8278).
edge(8278, 8279).
edge(8279, 8280).
edge(8280, 8281).
edge(8281, 8282).
edge(8282, 8283).
edge(8283, 8284).
edge(8284, 8285).
edge(8285, 8286).
edge(8286, 8287).
edge(8287, 8288).
edge(8288, 8289).
edge(8289, 8290).
edge(8290, 8291).
edge(8291, 8292).
edge(8292, 8293).
edge(8293, 8294).
edge(8294, 8295).
edge(8295, 8296).
edge(8296, 8297).
edge(8297, 8298).
edge(8298, 8299).
edge(8299, 8300).
edge(8300, 8301).
edge(8301, 8302).
edge(8302, 8303).
edge(8303, 8304).
edge(8304, 8305).
edge(8305, 8306).
edge(8306, 8307).
edge(8307, 8308).
edge(8308, 8309).
edge(8309, 8310).
edge(8310, 8311).
edge(8311, 8312).
edge(8312, 8313).
edge(8313, 8314).
edge(8314, 8315).
edge(8315, 8316).
edge(8316, 8317).
edge(8317, 8318).
edge(8318, 8319).
edge(8319, 8320).
edge(8320, 8321).
edge(8321, 8322).
edge(8322, 8323).
edge(8323, 8324).
edge(8324, 8325).
edge(8325, 8326).
edge(8326, 8327).
edge(8327, 8328).
edge(8328, 8329).
edge(8329, 8330).
edge(8330, 8331).
edge(8331, 8332).
edge(8332, 8333).
edge(8333, 8334).
edge(8334, 8335).
edge(8335, 8336).
edge(8336, 8337).
edge(8337, 8338).
edge(8338, 8339).
edge(8339, 8340).
edge(8340, 8341).
edge(8341, 8342).
edge(8342, 8343).
edge(8343, 8344).
edge(8344, 8345).
edge(8345, 8346).
edge(8346, 8347).
edge(8347, 8348).
edge(8348, 8349).
edge(8349, 8350).
edge(8350, 8351).
edge(8351, 8352).
edge(8352, 8353).
edge(8353, 8354).
edge(8354, 8355).
edge(8355, 8356).
edge(8356, 8357).
edge(8357, 8358).
edge(8358, 8359).
edge(8359, 8360).
edge(8360, 8361).
edge(8361, 8362).
edge(8362, 8363).
edge(8363, 8364).
edge(8364, 8365).
edge(8365, 8366).
edge(8366, 8367).
edge(8367, 8368).
edge(8368, 8369).
edge(8369, 8370).
edge(8370, 8371).
edge(8371, 8372).
edge(8372, 8373).
edge(8373, 8374).
edge(8374, 8375).
edge(8375, 8376).
edge(8376, 8377).
edge(8377, 8378).
edge(8378, 8379).
edge(8379, 8380).
edge(8380, 8381).
edge(8381, 8382).
edge(8382, 8383).
edge(8383, 8384).
edge(8384, 8385).
edge(8385, 8386).
edge(8386, 8387).
edge(8387, 8388).
edge(8388, 8389).
edge(8389, 8390).
edge(8390, 8391).
edge(8391, 8392).
edge(8392, 8393).
edge(8393, 8394).
edge(8394, 8395).
edge(8395, 8396).
edge(8396, 8397).
edge(8397, 8398).
edge(8398, 8399).
edge(8399, 8400).
edge(8400, 8401).
edge(8401, 8402).
edge(8402, 8403).
edge(8403, 8404).
edge(8404, 8405).
edge(8405, 8406).
edge(8406, 8407).
edge(8407, 8408).
edge(8408, 8409).
edge(8409, 8410).
edge(8410, 8411).
edge(8411, 8412).
edge(8412, 8413).
edge(8413, 8414).
edge(8414, 8415).
edge(8415, 8416).
edge(8416, 8417).
edge(8417, 8418).
edge(8418, 8419).
edge(8419, 8420).
edge(8420, 8421).
edge(8421, 8422).
edge(8422, 8423).
edge(8423, 8424).
edge(8424, 8425).
edge(8425, 8426).
edge(8426, 8427).
edge(8427, 8428).
edge(8428, 8429).
edge(8429, 8430).
edge(8430, 8431).
edge(8431, 8432).
edge(8432, 8433).
edge(8433, 8434).
edge(8434, 8435).
edge(8435, 8436).
edge(8436, 8437).
edge(8437, 8438).
edge(8438, 8439).
edge(8439, 8440).
edge(8440, 8441).
edge(8441, 8442).
edge(8442, 8443).
edge(8443, 8444).
edge(8444, 8445).
edge(8445, 8446).
edge(8446, 8447).
edge(8447, 8448).
edge(8448, 8449).
edge(8449, 8450).
edge(8450, 8451).
edge(8451, 8452).
edge(8452, 8453).
edge(8453, 8454).
edge(8454, 8455).
edge(8455, 8456).
edge(8456, 8457).
edge(8457, 8458).
edge(8458, 8459).
edge(8459, 8460).
edge(8460, 8461).
edge(8461, 8462).
edge(8462, 8463).
edge(8463, 8464).
edge(8464, 8465).
edge(8465, 8466).
edge(8466, 8467).
edge(8467, 8468).
edge(8468, 8469).
edge(8469, 8470).
edge(8470, 8471).
edge(8471, 8472).
edge(8472, 8473).
edge(8473, 8474).
edge(8474, 8475).
edge(8475, 8476).
edge(8476, 8477).
edge(8477, 8478).
edge(8478, 8479).
edge(8479, 8480).
edge(8480, 8481).
edge(8481, 8482).
edge(8482, 8483).
edge(8483, 8484).
edge(8484, 8485).
edge(8485, 8486).
edge(8486, 8487).
edge(8487, 8488).
edge(8488, 8489).
edge(8489, 8490).
edge(8490, 8491).
edge(8491, 8492).
edge(8492, 8493).
edge(8493, 8494).
edge(8494, 8495).
edge(8495, 8496).
edge(8496, 8497).
edge(8497, 8498).
edge(8498, 8499).
edge(8499, 8500).
edge(8500, 8501).
edge(8501, 8502).
edge(8502, 8503).
edge(8503, 8504).
edge(8504, 8505).
edge(8505, 8506).
edge(8506, 8507).
edge(8507, 8508).
edge(8508, 8509).
edge(8509, 8510).
edge(8510, 8511).
edge(8511, 8512).
edge(8512, 8513).
edge(8513, 8514).
edge(8514, 8515).
edge(8515, 8516).
edge(8516, 8517).
edge(8517, 8518).
edge(8518, 8519).
edge(8519, 8520).
edge(8520, 8521).
edge(8521, 8522).
edge(8522, 8523).
edge(8523, 8524).
edge(8524, 8525).
edge(8525, 8526).
edge(8526, 8527).
edge(8527, 8528).
edge(8528, 8529).
edge(8529, 8530).
edge(8530, 8531).
edge(8531, 8532).
edge(8532, 8533).
edge(8533, 8534).
edge(8534, 8535).
edge(8535, 8536).
edge(8536, 8537).
edge(8537, 8538).
edge(8538, 8539).
edge(8539, 8540).
edge(8540, 8541).
edge(8541, 8542).
edge(8542, 8543).
edge(8543, 8544).
edge(8544, 8545).
edge(8545, 8546).
edge(8546, 8547).
edge(8547, 8548).
edge(8548, 8549).
edge(8549, 8550).
edge(8550, 8551).
edge(8551, 8552).
edge(8552, 8553).
edge(8553, 8554).
edge(8554, 8555).
edge(8555, 8556).
edge(8556, 8557).
edge(8557, 8558).
edge(8558, 8559).
edge(8559, 8560).
edge(8560, 8561).
edge(8561, 8562).
edge(8562, 8563).
edge(8563, 8564).
edge(8564, 8565).
edge(8565, 8566).
edge(8566, 8567).
edge(8567, 8568).
edge(8568, 8569).
edge(8569, 8570).
edge(8570, 8571).
edge(8571, 8572).
edge(8572, 8573).
edge(8573, 8574).
edge(8574, 8575).
edge(8575, 8576).
edge(8576, 8577).
edge(8577, 8578).
edge(8578, 8579).
edge(8579, 8580).
edge(8580, 8581).
edge(8581, 8582).
edge(8582, 8583).
edge(8583, 8584).
edge(8584, 8585).
edge(8585, 8586).
edge(8586, 8587).
edge(8587, 8588).
edge(8588, 8589).
edge(8589, 8590).
edge(8590, 8591).
edge(8591, 8592).
edge(8592, 8593).
edge(8593, 8594).
edge(8594, 8595).
edge(8595, 8596).
edge(8596, 8597).
edge(8597, 8598).
edge(8598, 8599).
edge(8599, 8600).
edge(8600, 8601).
edge(8601, 8602).
edge(8602, 8603).
edge(8603, 8604).
edge(8604, 8605).
edge(8605, 8606).
edge(8606, 8607).
edge(8607, 8608).
edge(8608, 8609).
edge(8609, 8610).
edge(8610, 8611).
edge(8611, 8612).
edge(8612, 8613).
edge(8613, 8614).
edge(8614, 8615).
edge(8615, 8616).
edge(8616, 8617).
edge(8617, 8618).
edge(8618, 8619).
edge(8619, 8620).
edge(8620, 8621).
edge(8621, 8622).
edge(8622, 8623).
edge(8623, 8624).
edge(8624, 8625).
edge(8625, 8626).
edge(8626, 8627).
edge(8627, 8628).
edge(8628, 8629).
edge(8629, 8630).
edge(8630, 8631).
edge(8631, 8632).
edge(8632, 8633).
edge(8633, 8634).
edge(8634, 8635).
edge(8635, 8636).
edge(8636, 8637).
edge(8637, 8638).
edge(8638, 8639).
edge(8639, 8640).
edge(8640, 8641).
edge(8641, 8642).
edge(8642, 8643).
edge(8643, 8644).
edge(8644, 8645).
edge(8645, 8646).
edge(8646, 8647).
edge(8647, 8648).
edge(8648, 8649).
edge(8649, 8650).
edge(8650, 8651).
edge(8651, 8652).
edge(8652, 8653).
edge(8653, 8654).
edge(8654, 8655).
edge(8655, 8656).
edge(8656, 8657).
edge(8657, 8658).
edge(8658, 8659).
edge(8659, 8660).
edge(8660, 8661).
edge(8661, 8662).
edge(8662, 8663).
edge(8663, 8664).
edge(8664, 8665).
edge(8665, 8666).
edge(8666, 8667).
edge(8667, 8668).
edge(8668, 8669).
edge(8669, 8670).
edge(8670, 8671).
edge(8671, 8672).
edge(8672, 8673).
edge(8673, 8674).
edge(8674, 8675).
edge(8675, 8676).
edge(8676, 8677).
edge(8677, 8678).
edge(8678, 8679).
edge(8679, 8680).
edge(8680, 8681).
edge(8681, 8682).
edge(8682, 8683).
edge(8683, 8684).
edge(8684, 8685).
edge(8685, 8686).
edge(8686, 8687).
edge(8687, 8688).
edge(8688, 8689).
edge(8689, 8690).
edge(8690, 8691).
edge(8691, 8692).
edge(8692, 8693).
edge(8693, 8694).
edge(8694, 8695).
edge(8695, 8696).
edge(8696, 8697).
edge(8697, 8698).
edge(8698, 8699).
edge(8699, 8700).
edge(8700, 8701).
edge(8701, 8702).
edge(8702, 8703).
edge(8703, 8704).
edge(8704, 8705).
edge(8705, 8706).
edge(8706, 8707).
edge(8707, 8708).
edge(8708, 8709).
edge(8709, 8710).
edge(8710, 8711).
edge(8711, 8712).
edge(8712, 8713).
edge(8713, 8714).
edge(8714, 8715).
edge(8715, 8716).
edge(8716, 8717).
edge(8717, 8718).
edge(8718, 8719).
edge(8719, 8720).
edge(8720, 8721).
edge(8721, 8722).
edge(8722, 8723).
edge(8723, 8724).
edge(8724, 8725).
edge(8725, 8726).
edge(8726, 8727).
edge(8727, 8728).
edge(8728, 8729).
edge(8729, 8730).
edge(8730, 8731).
edge(8731, 8732).
edge(8732, 8733).
edge(8733, 8734).
edge(8734, 8735).
edge(8735, 8736).
edge(8736, 8737).
edge(8737, 8738).
edge(8738, 8739).
edge(8739, 8740).
edge(8740, 8741).
edge(8741, 8742).
edge(8742, 8743).
edge(8743, 8744).
edge(8744, 8745).
edge(8745, 8746).
edge(8746, 8747).
edge(8747, 8748).
edge(8748, 8749).
edge(8749, 8750).
edge(8750, 8751).
edge(8751, 8752).
edge(8752, 8753).
edge(8753, 8754).
edge(8754, 8755).
edge(8755, 8756).
edge(8756, 8757).
edge(8757, 8758).
edge(8758, 8759).
edge(8759, 8760).
edge(8760, 8761).
edge(8761, 8762).
edge(8762, 8763).
edge(8763, 8764).
edge(8764, 8765).
edge(8765, 8766).
edge(8766, 8767).
edge(8767, 8768).
edge(8768, 8769).
edge(8769, 8770).
edge(8770, 8771).
edge(8771, 8772).
edge(8772, 8773).
edge(8773, 8774).
edge(8774, 8775).
edge(8775, 8776).
edge(8776, 8777).
edge(8777, 8778).
edge(8778, 8779).
edge(8779, 8780).
edge(8780, 8781).
edge(8781, 8782).
edge(8782, 8783).
edge(8783, 8784).
edge(8784, 8785).
edge(8785, 8786).
edge(8786, 8787).
edge(8787, 8788).
edge(8788, 8789).
edge(8789, 8790).
edge(8790, 8791).
edge(8791, 8792).
edge(8792, 8793).
edge(8793, 8794).
edge(8794, 8795).
edge(8795, 8796).
edge(8796, 8797).
edge(8797, 8798).
edge(8798, 8799).
edge(8799, 8800).
edge(8800, 8801).
edge(8801, 8802).
edge(8802, 8803).
edge(8803, 8804).
edge(8804, 8805).
edge(8805, 8806).
edge(8806, 8807).
edge(8807, 8808).
edge(8808, 8809).
edge(8809, 8810).
edge(8810, 8811).
edge(8811, 8812).
edge(8812, 8813).
edge(8813, 8814).
edge(8814, 8815).
edge(8815, 8816).
edge(8816, 8817).
edge(8817, 8818).
edge(8818, 8819).
edge(8819, 8820).
edge(8820, 8821).
edge(8821, 8822).
edge(8822, 8823).
edge(8823, 8824).
edge(8824, 8825).
edge(8825, 8826).
edge(8826, 8827).
edge(8827, 8828).
edge(8828, 8829).
edge(8829, 8830).
edge(8830, 8831).
edge(8831, 8832).
edge(8832, 8833).
edge(8833, 8834).
edge(8834, 8835).
edge(8835, 8836).
edge(8836, 8837).
edge(8837, 8838).
edge(8838, 8839).
edge(8839, 8840).
edge(8840, 8841).
edge(8841, 8842).
edge(8842, 8843).
edge(8843, 8844).
edge(8844, 8845).
edge(8845, 8846).
edge(8846, 8847).
edge(8847, 8848).
edge(8848, 8849).
edge(8849, 8850).
edge(8850, 8851).
edge(8851, 8852).
edge(8852, 8853).
edge(8853, 8854).
edge(8854, 8855).
edge(8855, 8856).
edge(8856, 8857).
edge(8857, 8858).
edge(8858, 8859).
edge(8859, 8860).
edge(8860, 8861).
edge(8861, 8862).
edge(8862, 8863).
edge(8863, 8864).
edge(8864, 8865).
edge(8865, 8866).
edge(8866, 8867).
edge(8867, 8868).
edge(8868, 8869).
edge(8869, 8870).
edge(8870, 8871).
edge(8871, 8872).
edge(8872, 8873).
edge(8873, 8874).
edge(8874, 8875).
edge(8875, 8876).
edge(8876, 8877).
edge(8877, 8878).
edge(8878, 8879).
edge(8879, 8880).
edge(8880, 8881).
edge(8881, 8882).
edge(8882, 8883).
edge(8883, 8884).
edge(8884, 8885).
edge(8885, 8886).
edge(8886, 8887).
edge(8887, 8888).
edge(8888, 8889).
edge(8889, 8890).
edge(8890, 8891).
edge(8891, 8892).
edge(8892, 8893).
edge(8893, 8894).
edge(8894, 8895).
edge(8895, 8896).
edge(8896, 8897).
edge(8897, 8898).
edge(8898, 8899).
edge(8899, 8900).
edge(8900, 8901).
edge(8901, 8902).
edge(8902, 8903).
edge(8903, 8904).
edge(8904, 8905).
edge(8905, 8906).
edge(8906, 8907).
edge(8907, 8908).
edge(8908, 8909).
edge(8909, 8910).
edge(8910, 8911).
edge(8911, 8912).
edge(8912, 8913).
edge(8913, 8914).
edge(8914, 8915).
edge(8915, 8916).
edge(8916, 8917).
edge(8917, 8918).
edge(8918, 8919).
edge(8919, 8920).
edge(8920, 8921).
edge(8921, 8922).
edge(8922, 8923).
edge(8923, 8924).
edge(8924, 8925).
edge(8925, 8926).
edge(8926, 8927).
edge(8927, 8928).
edge(8928, 8929).
edge(8929, 8930).
edge(8930, 8931).
edge(8931, 8932).
edge(8932, 8933).
edge(8933, 8934).
edge(8934, 8935).
edge(8935, 8936).
edge(8936, 8937).
edge(8937, 8938).
edge(8938, 8939).
edge(8939, 8940).
edge(8940, 8941).
edge(8941, 8942).
edge(8942, 8943).
edge(8943, 8944).
edge(8944, 8945).
edge(8945, 8946).
edge(8946, 8947).
edge(8947, 8948).
edge(8948, 8949).
edge(8949, 8950).
edge(8950, 8951).
edge(8951, 8952).
edge(8952, 8953).
edge(8953, 8954).
edge(8954, 8955).
edge(8955, 8956).
edge(8956, 8957).
edge(8957, 8958).
edge(8958, 8959).
edge(8959, 8960).
edge(8960, 8961).
edge(8961, 8962).
edge(8962, 8963).
edge(8963, 8964).
edge(8964, 8965).
edge(8965, 8966).
edge(8966, 8967).
edge(8967, 8968).
edge(8968, 8969).
edge(8969, 8970).
edge(8970, 8971).
edge(8971, 8972).
edge(8972, 8973).
edge(8973, 8974).
edge(8974, 8975).
edge(8975, 8976).
edge(8976, 8977).
edge(8977, 8978).
edge(8978, 8979).
edge(8979, 8980).
edge(8980, 8981).
edge(8981, 8982).
edge(8982, 8983).
edge(8983, 8984).
edge(8984, 8985).
edge(8985, 8986).
edge(8986, 8987).
edge(8987, 8988).
edge(8988, 8989).
edge(8989, 8990).
edge(8990, 8991).
edge(8991, 8992).
edge(8992, 8993).
edge(8993, 8994).
edge(8994, 8995).
edge(8995, 8996).
edge(8996, 8997).
edge(8997, 8998).
edge(8998, 8999).
edge(8999, 9000).
edge(9000, 9001).
edge(9001, 9002).
edge(9002, 9003).
edge(9003, 9004).
edge(9004, 9005).
edge(9005, 9006).
edge(9006, 9007).
edge(9007, 9008).
edge(9008, 9009).
edge(9009, 9010).
edge(9010, 9011).
edge(9011, 9012).
edge(9012, 9013).
edge(9013, 9014).
edge(9014, 9015).
edge(9015, 9016).
edge(9016, 9017).
edge(9017, 9018).
edge(9018, 9019).
edge(9019, 9020).
edge(9020, 9021).
edge(9021, 9022).
edge(9022, 9023).
edge(9023, 9024).
edge(9024, 9025).
edge(9025, 9026).
edge(9026, 9027).
edge(9027, 9028).
edge(9028, 9029).
edge(9029, 9030).
edge(9030, 9031).
edge(9031, 9032).
edge(9032, 9033).
edge(9033, 9034).
edge(9034, 9035).
edge(9035, 9036).
edge(9036, 9037).
edge(9037, 9038).
edge(9038, 9039).
edge(9039, 9040).
edge(9040, 9041).
edge(9041, 9042).
edge(9042, 9043).
edge(9043, 9044).
edge(9044, 9045).
edge(9045, 9046).
edge(9046, 9047).
edge(9047, 9048).
edge(9048, 9049).
edge(9049, 9050).
edge(9050, 9051).
edge(9051, 9052).
edge(9052, 9053).
edge(9053, 9054).
edge(9054, 9055).
edge(9055, 9056).
edge(9056, 9057).
edge(9057, 9058).
edge(9058, 9059).
edge(9059, 9060).
edge(9060, 9061).
edge(9061, 9062).
edge(9062, 9063).
edge(9063, 9064).
edge(9064, 9065).
edge(9065, 9066).
edge(9066, 9067).
edge(9067, 9068).
edge(9068, 9069).
edge(9069, 9070).
edge(9070, 9071).
edge(9071, 9072).
edge(9072, 9073).
edge(9073, 9074).
edge(9074, 9075).
edge(9075, 9076).
edge(9076, 9077).
edge(9077, 9078).
edge(9078, 9079).
edge(9079, 9080).
edge(9080, 9081).
edge(9081, 9082).
edge(9082, 9083).
edge(9083, 9084).
edge(9084, 9085).
edge(9085, 9086).
edge(9086, 9087).
edge(9087, 9088).
edge(9088, 9089).
edge(9089, 9090).
edge(9090, 9091).
edge(9091, 9092).
edge(9092, 9093).
edge(9093, 9094).
edge(9094, 9095).
edge(9095, 9096).
edge(9096, 9097).
edge(9097, 9098).
edge(9098, 9099).
edge(9099, 9100).
edge(9100, 9101).
edge(9101, 9102).
edge(9102, 9103).
edge(9103, 9104).
edge(9104, 9105).
edge(9105, 9106).
edge(9106, 9107).
edge(9107, 9108).
edge(9108, 9109).
edge(9109, 9110).
edge(9110, 9111).
edge(9111, 9112).
edge(9112, 9113).
edge(9113, 9114).
edge(9114, 9115).
edge(9115, 9116).
edge(9116, 9117).
edge(9117, 9118).
edge(9118, 9119).
edge(9119, 9120).
edge(9120, 9121).
edge(9121, 9122).
edge(9122, 9123).
edge(9123, 9124).
edge(9124, 9125).
edge(9125, 9126).
edge(9126, 9127).
edge(9127, 9128).
edge(9128, 9129).
edge(9129, 9130).
edge(9130, 9131).
edge(9131, 9132).
edge(9132, 9133).
edge(9133, 9134).
edge(9134, 9135).
edge(9135, 9136).
edge(9136, 9137).
edge(9137, 9138).
edge(9138, 9139).
edge(9139, 9140).
edge(9140, 9141).
edge(9141, 9142).
edge(9142, 9143).
edge(9143, 9144).
edge(9144, 9145).
edge(9145, 9146).
edge(9146, 9147).
edge(9147, 9148).
edge(9148, 9149).
edge(9149, 9150).
edge(9150, 9151).
edge(9151, 9152).
edge(9152, 9153).
edge(9153, 9154).
edge(9154, 9155).
edge(9155, 9156).
edge(9156, 9157).
edge(9157, 9158).
edge(9158, 9159).
edge(9159, 9160).
edge(9160, 9161).
edge(9161, 9162).
edge(9162, 9163).
edge(9163, 9164).
edge(9164, 9165).
edge(9165, 9166).
edge(9166, 9167).
edge(9167, 9168).
edge(9168, 9169).
edge(9169, 9170).
edge(9170, 9171).
edge(9171, 9172).
edge(9172, 9173).
edge(9173, 9174).
edge(9174, 9175).
edge(9175, 9176).
edge(9176, 9177).
edge(9177, 9178).
edge(9178, 9179).
edge(9179, 9180).
edge(9180, 9181).
edge(9181, 9182).
edge(9182, 9183).
edge(9183, 9184).
edge(9184, 9185).
edge(9185, 9186).
edge(9186, 9187).
edge(9187, 9188).
edge(9188, 9189).
edge(9189, 9190).
edge(9190, 9191).
edge(9191, 9192).
edge(9192, 9193).
edge(9193, 9194).
edge(9194, 9195).
edge(9195, 9196).
edge(9196, 9197).
edge(9197, 9198).
edge(9198, 9199).
edge(9199, 9200).
edge(9200, 9201).
edge(9201, 9202).
edge(9202, 9203).
edge(9203, 9204).
edge(9204, 9205).
edge(9205, 9206).
edge(9206, 9207).
edge(9207, 9208).
edge(9208, 9209).
edge(9209, 9210).
edge(9210, 9211).
edge(9211, 9212).
edge(9212, 9213).
edge(9213, 9214).
edge(9214, 9215).
edge(9215, 9216).
edge(9216, 9217).
edge(9217, 9218).
edge(9218, 9219).
edge(9219, 9220).
edge(9220, 9221).
edge(9221, 9222).
edge(9222, 9223).
edge(9223, 9224).
edge(9224, 9225).
edge(9225, 9226).
edge(9226, 9227).
edge(9227, 9228).
edge(9228, 9229).
edge(9229, 9230).
edge(9230, 9231).
edge(9231, 9232).
edge(9232, 9233).
edge(9233, 9234).
edge(9234, 9235).
edge(9235, 9236).
edge(9236, 9237).
edge(9237, 9238).
edge(9238, 9239).
edge(9239, 9240).
edge(9240, 9241).
edge(9241, 9242).
edge(9242, 9243).
edge(9243, 9244).
edge(9244, 9245).
edge(9245, 9246).
edge(9246, 9247).
edge(9247, 9248).
edge(9248, 9249).
edge(9249, 9250).
edge(9250, 9251).
edge(9251, 9252).
edge(9252, 9253).
edge(9253, 9254).
edge(9254, 9255).
edge(9255, 9256).
edge(9256, 9257).
edge(9257, 9258).
edge(9258, 9259).
edge(9259, 9260).
edge(9260, 9261).
edge(9261, 9262).
edge(9262, 9263).
edge(9263, 9264).
edge(9264, 9265).
edge(9265, 9266).
edge(9266, 9267).
edge(9267, 9268).
edge(9268, 9269).
edge(9269, 9270).
edge(9270, 9271).
edge(9271, 9272).
edge(9272, 9273).
edge(9273, 9274).
edge(9274, 9275).
edge(9275, 9276).
edge(9276, 9277).
edge(9277, 9278).
edge(9278, 9279).
edge(9279, 9280).
edge(9280, 9281).
edge(9281, 9282).
edge(9282, 9283).
edge(9283, 9284).
edge(9284, 9285).
edge(9285, 9286).
edge(9286, 9287).
edge(9287, 9288).
edge(9288, 9289).
edge(9289, 9290).
edge(9290, 9291).
edge(9291, 9292).
edge(9292, 9293).
edge(9293, 9294).
edge(9294, 9295).
edge(9295, 9296).
edge(9296, 9297).
edge(9297, 9298).
edge(9298, 9299).
edge(9299, 9300).
edge(9300, 9301).
edge(9301, 9302).
edge(9302, 9303).
edge(9303, 9304).
edge(9304, 9305).
edge(9305, 9306).
edge(9306, 9307).
edge(9307, 9308).
edge(9308, 9309).
edge(9309, 9310).
edge(9310, 9311).
edge(9311, 9312).
edge(9312, 9313).
edge(9313, 9314).
edge(9314, 9315).
edge(9315, 9316).
edge(9316, 9317).
edge(9317, 9318).
edge(9318, 9319).
edge(9319, 9320).
edge(9320, 9321).
edge(9321, 9322).
edge(9322, 9323).
edge(9323, 9324).
edge(9324, 9325).
edge(9325, 9326).
edge(9326, 9327).
edge(9327, 9328).
edge(9328, 9329).
edge(9329, 9330).
edge(9330, 9331).
edge(9331, 9332).
edge(9332, 9333).
edge(9333, 9334).
edge(9334, 9335).
edge(9335, 9336).
edge(9336, 9337).
edge(9337, 9338).
edge(9338, 9339).
edge(9339, 9340).
edge(9340, 9341).
edge(9341, 9342).
edge(9342, 9343).
edge(9343, 9344).
edge(9344, 9345).
edge(9345, 9346).
edge(9346, 9347).
edge(9347, 9348).
edge(9348, 9349).
edge(9349, 9350).
edge(9350, 9351).
edge(9351, 9352).
edge(9352, 9353).
edge(9353, 9354).
edge(9354, 9355).
edge(9355, 9356).
edge(9356, 9357).
edge(9357, 9358).
edge(9358, 9359).
edge(9359, 9360).
edge(9360, 9361).
edge(9361, 9362).
edge(9362, 9363).
edge(9363, 9364).
edge(9364, 9365).
edge(9365, 9366).
edge(9366, 9367).
edge(9367, 9368).
edge(9368, 9369).
edge(9369, 9370).
edge(9370, 9371).
edge(9371, 9372).
edge(9372, 9373).
edge(9373, 9374).
edge(9374, 9375).
edge(9375, 9376).
edge(9376, 9377).
edge(9377, 9378).
edge(9378, 9379).
edge(9379, 9380).
edge(9380, 9381).
edge(9381, 9382).
edge(9382, 9383).
edge(9383, 9384).
edge(9384, 9385).
edge(9385, 9386).
edge(9386, 9387).
edge(9387, 9388).
edge(9388, 9389).
edge(9389, 9390).
edge(9390, 9391).
edge(9391, 9392).
edge(9392, 9393).
edge(9393, 9394).
edge(9394, 9395).
edge(9395, 9396).
edge(9396, 9397).
edge(9397, 9398).
edge(9398, 9399).
edge(9399, 9400).
edge(9400, 9401).
edge(9401, 9402).
edge(9402, 9403).
edge(9403, 9404).
edge(9404, 9405).
edge(9405, 9406).
edge(9406, 9407).
edge(9407, 9408).
edge(9408, 9409).
edge(9409, 9410).
edge(9410, 9411).
edge(9411, 9412).
edge(9412, 9413).
edge(9413, 9414).
edge(9414, 9415).
edge(9415, 9416).
edge(9416, 9417).
edge(9417, 9418).
edge(9418, 9419).
edge(9419, 9420).
edge(9420, 9421).
edge(9421, 9422).
edge(9422, 9423).
edge(9423, 9424).
edge(9424, 9425).
edge(9425, 9426).
edge(9426, 9427).
edge(9427, 9428).
edge(9428, 9429).
edge(9429, 9430).
edge(9430, 9431).
edge(9431, 9432).
edge(9432, 9433).
edge(9433, 9434).
edge(9434, 9435).
edge(9435, 9436).
edge(9436, 9437).
edge(9437, 9438).
edge(9438, 9439).
edge(9439, 9440).
edge(9440, 9441).
edge(9441, 9442).
edge(9442, 9443).
edge(9443, 9444).
edge(9444, 9445).
edge(9445, 9446).
edge(9446, 9447).
edge(9447, 9448).
edge(9448, 9449).
edge(9449, 9450).
edge(9450, 9451).
edge(9451, 9452).
edge(9452, 9453).
edge(9453, 9454).
edge(9454, 9455).
edge(9455, 9456).
edge(9456, 9457).
edge(9457, 9458).
edge(9458, 9459).
edge(9459, 9460).
edge(9460, 9461).
edge(9461, 9462).
edge(9462, 9463).
edge(9463, 9464).
edge(9464, 9465).
edge(9465, 9466).
edge(9466, 9467).
edge(9467, 9468).
edge(9468, 9469).
edge(9469, 9470).
edge(9470, 9471).
edge(9471, 9472).
edge(9472, 9473).
edge(9473, 9474).
edge(9474, 9475).
edge(9475, 9476).
edge(9476, 9477).
edge(9477, 9478).
edge(9478, 9479).
edge(9479, 9480).
edge(9480, 9481).
edge(9481, 9482).
edge(9482, 9483).
edge(9483, 9484).
edge(9484, 9485).
edge(9485, 9486).
edge(9486, 9487).
edge(9487, 9488).
edge(9488, 9489).
edge(9489, 9490).
edge(9490, 9491).
edge(9491, 9492).
edge(9492, 9493).
edge(9493, 9494).
edge(9494, 9495).
edge(9495, 9496).
edge(9496, 9497).
edge(9497, 9498).
edge(9498, 9499).
edge(9499, 9500).
edge(9500, 9501).
edge(9501, 9502).
edge(9502, 9503).
edge(9503, 9504).
edge(9504, 9505).
edge(9505, 9506).
edge(9506, 9507).
edge(9507, 9508).
edge(9508, 9509).
edge(9509, 9510).
edge(9510, 9511).
edge(9511, 9512).
edge(9512, 9513).
edge(9513, 9514).
edge(9514, 9515).
edge(9515, 9516).
edge(9516, 9517).
edge(9517, 9518).
edge(9518, 9519).
edge(9519, 9520).
edge(9520, 9521).
edge(9521, 9522).
edge(9522, 9523).
edge(9523, 9524).
edge(9524, 9525).
edge(9525, 9526).
edge(9526, 9527).
edge(9527, 9528).
edge(9528, 9529).
edge(9529, 9530).
edge(9530, 9531).
edge(9531, 9532).
edge(9532, 9533).
edge(9533, 9534).
edge(9534, 9535).
edge(9535, 9536).
edge(9536, 9537).
edge(9537, 9538).
edge(9538, 9539).
edge(9539, 9540).
edge(9540, 9541).
edge(9541, 9542).
edge(9542, 9543).
edge(9543, 9544).
edge(9544, 9545).
edge(9545, 9546).
edge(9546, 9547).
edge(9547, 9548).
edge(9548, 9549).
edge(9549, 9550).
edge(9550, 9551).
edge(9551, 9552).
edge(9552, 9553).
edge(9553, 9554).
edge(9554, 9555).
edge(9555, 9556).
edge(9556, 9557).
edge(9557, 9558).
edge(9558, 9559).
edge(9559, 9560).
edge(9560, 9561).
edge(9561, 9562).
edge(9562, 9563).
edge(9563, 9564).
edge(9564, 9565).
edge(9565, 9566).
edge(9566, 9567).
edge(9567, 9568).
edge(9568, 9569).
edge(9569, 9570).
edge(9570, 9571).
edge(9571, 9572).
edge(9572, 9573).
edge(9573, 9574).
edge(9574, 9575).
edge(9575, 9576).
edge(9576, 9577).
edge(9577, 9578).
edge(9578, 9579).
edge(9579, 9580).
edge(9580, 9581).
edge(9581, 9582).
edge(9582, 9583).
edge(9583, 9584).
edge(9584, 9585).
edge(9585, 9586).
edge(9586, 9587).
edge(9587, 9588).
edge(9588, 9589).
edge(9589, 9590).
edge(9590, 9591).
edge(9591, 9592).
edge(9592, 9593).
edge(9593, 9594).
edge(9594, 9595).
edge(9595, 9596).
edge(9596, 9597).
edge(9597, 9598).
edge(9598, 9599).
edge(9599, 9600).
edge(9600, 9601).
edge(9601, 9602).
edge(9602, 9603).
edge(9603, 9604).
edge(9604, 9605).
edge(9605, 9606).
edge(9606, 9607).
edge(9607, 9608).
edge(9608, 9609).
edge(9609, 9610).
edge(9610, 9611).
edge(9611, 9612).
edge(9612, 9613).
edge(9613, 9614).
edge(9614, 9615).
edge(9615, 9616).
edge(9616, 9617).
edge(9617, 9618).
edge(9618, 9619).
edge(9619, 9620).
edge(9620, 9621).
edge(9621, 9622).
edge(9622, 9623).
edge(9623, 9624).
edge(9624, 9625).
edge(9625, 9626).
edge(9626, 9627).
edge(9627, 9628).
edge(9628, 9629).
edge(9629, 9630).
edge(9630, 9631).
edge(9631, 9632).
edge(9632, 9633).
edge(9633, 9634).
edge(9634, 9635).
edge(9635, 9636).
edge(9636, 9637).
edge(9637, 9638).
edge(9638, 9639).
edge(9639, 9640).
edge(9640, 9641).
edge(9641, 9642).
edge(9642, 9643).
edge(9643, 9644).
edge(9644, 9645).
edge(9645, 9646).
edge(9646, 9647).
edge(9647, 9648).
edge(9648, 9649).
edge(9649, 9650).
edge(9650, 9651).
edge(9651, 9652).
edge(9652, 9653).
edge(9653, 9654).
edge(9654, 9655).
edge(9655, 9656).
edge(9656, 9657).
edge(9657, 9658).
edge(9658, 9659).
edge(9659, 9660).
edge(9660, 9661).
edge(9661, 9662).
edge(9662, 9663).
edge(9663, 9664).
edge(9664, 9665).
edge(9665, 9666).
edge(9666, 9667).
edge(9667, 9668).
edge(9668, 9669).
edge(9669, 9670).
edge(9670, 9671).
edge(9671, 9672).
edge(9672, 9673).
edge(9673, 9674).
edge(9674, 9675).
edge(9675, 9676).
edge(9676, 9677).
edge(9677, 9678).
edge(9678, 9679).
edge(9679, 9680).
edge(9680, 9681).
edge(9681, 9682).
edge(9682, 9683).
edge(9683, 9684).
edge(9684, 9685).
edge(9685, 9686).
edge(9686, 9687).
edge(9687, 9688).
edge(9688, 9689).
edge(9689, 9690).
edge(9690, 9691).
edge(9691, 9692).
edge(9692, 9693).
edge(9693, 9694).
edge(9694, 9695).
edge(9695, 9696).
edge(9696, 9697).
edge(9697, 9698).
edge(9698, 9699).
edge(9699, 9700).
edge(9700, 9701).
edge(9701, 9702).
edge(9702, 9703).
edge(9703, 9704).
edge(9704, 9705).
edge(9705, 9706).
edge(9706, 9707).
edge(9707, 9708).
edge(9708, 9709).
edge(9709, 9710).
edge(9710, 9711).
edge(9711, 9712).
edge(9712, 9713).
edge(9713, 9714).
edge(9714, 9715).
edge(9715, 9716).
edge(9716, 9717).
edge(9717, 9718).
edge(9718, 9719).
edge(9719, 9720).
edge(9720, 9721).
edge(9721, 9722).
edge(9722, 9723).
edge(9723, 9724).
edge(9724, 9725).
edge(9725, 9726).
edge(9726, 9727).
edge(9727, 9728).
edge(9728, 9729).
edge(9729, 9730).
edge(9730, 9731).
edge(9731, 9732).
edge(9732, 9733).
edge(9733, 9734).
edge(9734, 9735).
edge(9735, 9736).
edge(9736, 9737).
edge(9737, 9738).
edge(9738, 9739).
edge(9739, 9740).
edge(9740, 9741).
edge(9741, 9742).
edge(9742, 9743).
edge(9743, 9744).
edge(9744, 9745).
edge(9745, 9746).
edge(9746, 9747).
edge(9747, 9748).
edge(9748, 9749).
edge(9749, 9750).
edge(9750, 9751).
edge(9751, 9752).
edge(9752, 9753).
edge(9753, 9754).
edge(9754, 9755).
edge(9755, 9756).
edge(9756, 9757).
edge(9757, 9758).
edge(9758, 9759).
edge(9759, 9760).
edge(9760, 9761).
edge(9761, 9762).
edge(9762, 9763).
edge(9763, 9764).
edge(9764, 9765).
edge(9765, 9766).
edge(9766, 9767).
edge(9767, 9768).
edge(9768, 9769).
edge(9769, 9770).
edge(9770, 9771).
edge(9771, 9772).
edge(9772, 9773).
edge(9773, 9774).
edge(9774, 9775).
edge(9775, 9776).
edge(9776, 9777).
edge(9777, 9778).
edge(9778, 9779).
edge(9779, 9780).
edge(9780, 9781).
edge(9781, 9782).
edge(9782, 9783).
edge(9783, 9784).
edge(9784, 9785).
edge(9785, 9786).
edge(9786, 9787).
edge(9787, 9788).
edge(9788, 9789).
edge(9789, 9790).
edge(9790, 9791).
edge(9791, 9792).
edge(9792, 9793).
edge(9793, 9794).
edge(9794, 9795).
edge(9795, 9796).
edge(9796, 9797).
edge(9797, 9798).
edge(9798, 9799).
edge(9799, 9800).
edge(9800, 9801).
edge(9801, 9802).
edge(9802, 9803).
edge(9803, 9804).
edge(9804, 9805).
edge(9805, 9806).
edge(9806, 9807).
edge(9807, 9808).
edge(9808, 9809).
edge(9809, 9810).
edge(9810, 9811).
edge(9811, 9812).
edge(9812, 9813).
edge(9813, 9814).
edge(9814, 9815).
edge(9815, 9816).
edge(9816, 9817).
edge(9817, 9818).
edge(9818, 9819).
edge(9819, 9820).
edge(9820, 9821).
edge(9821, 9822).
edge(9822, 9823).
edge(9823, 9824).
edge(9824, 9825).
edge(9825, 9826).
edge(9826, 9827).
edge(9827, 9828).
edge(9828, 9829).
edge(9829, 9830).
edge(9830, 9831).
edge(9831, 9832).
edge(9832, 9833).
edge(9833, 9834).
edge(9834, 9835).
edge(9835, 9836).
edge(9836, 9837).
edge(9837, 9838).
edge(9838, 9839).
edge(9839, 9840).
edge(9840, 9841).
edge(9841, 9842).
edge(9842, 9843).
edge(9843, 9844).
edge(9844, 9845).
edge(9845, 9846).
edge(9846, 9847).
edge(9847, 9848).
edge(9848, 9849).
edge(9849, 9850).
edge(9850, 9851).
edge(9851, 9852).
edge(9852, 9853).
edge(9853, 9854).
edge(9854, 9855).
edge(9855, 9856).
edge(9856, 9857).
edge(9857, 9858).
edge(9858, 9859).
edge(9859, 9860).
edge(9860, 9861).
edge(9861, 9862).
edge(9862, 9863).
edge(9863, 9864).
edge(9864, 9865).
edge(9865, 9866).
edge(9866, 9867).
edge(9867, 9868).
edge(9868, 9869).
edge(9869, 9870).
edge(9870, 9871).
edge(9871, 9872).
edge(9872, 9873).
edge(9873, 9874).
edge(9874, 9875).
edge(9875, 9876).
edge(9876, 9877).
edge(9877, 9878).
edge(9878, 9879).
edge(9879, 9880).
edge(9880, 9881).
edge(9881, 9882).
edge(9882, 9883).
edge(9883, 9884).
edge(9884, 9885).
edge(9885, 9886).
edge(9886, 9887).
edge(9887, 9888).
edge(9888, 9889).
edge(9889, 9890).
edge(9890, 9891).
edge(9891, 9892).
edge(9892, 9893).
edge(9893, 9894).
edge(9894, 9895).
edge(9895, 9896).
edge(9896, 9897).
edge(9897, 9898).
edge(9898, 9899).
edge(9899, 9900).
edge(9900, 9901).
edge(9901, 9902).
edge(9902, 9903).
edge(9903, 9904).
edge(9904, 9905).
edge(9905, 9906).
edge(9906, 9907).
edge(9907, 9908).
edge(9908, 9909).
edge(9909, 9910).
edge(9910, 9911).
edge(9911, 9912).
edge(9912, 9913).
edge(9913, 9914).
edge(9914, 9915).
edge(9915, 9916).
edge(9916, 9917).
edge(9917, 9918).
edge(9918, 9919).
edge(9919, 9920).
edge(9920, 9921).
edge(9921, 9922).
edge(9922, 9923).
edge(9923, 9924).
edge(9924, 9925).
edge(9925, 9926).
edge(9926, 9927).
edge(9927, 9928).
edge(9928, 9929).
edge(9929, 9930).
edge(9930, 9931).
edge(9931, 9932).
edge(9932, 9933).
edge(9933, 9934).
edge(9934, 9935).
edge(9935, 9936).
edge(9936, 9937).
edge(9937, 9938).
edge(9938, 9939).
edge(9939, 9940).
edge(9940, 9941).
edge(9941, 9942).
edge(9942, 9943).
edge(9943, 9944).
edge(9944, 9945).
edge(9945, 9946).
edge(9946, 9947).
edge(9947, 9948).
edge(9948, 9949).
edge(9949, 9950).
edge(9950, 9951).
edge(9951, 9952).
edge(9952, 9953).
edge(9953, 9954).
edge(9954, 9955).
edge(9955, 9956).
edge(9956, 9957).
edge(9957, 9958).
edge(9958, 9959).
edge(9959, 9960).
edge(9960, 9961).
edge(9961, 9962).
edge(9962, 9963).
edge(9963, 9964).
edge(9964, 9965).
edge(9965, 9966).
edge(9966, 9967).
edge(9967, 9968).
edge(9968, 9969).
edge(9969, 9970).
edge(9970, 9971).
edge(9971, 9972).
edge(9972, 9973).
edge(9973, 9974).
edge(9974, 9975).
edge(9975, 9976).
edge(9976, 9977).
edge(9977, 9978).
edge(9978, 9979).
edge(9979, 9980).
edge(9980, 9981).
edge(9981, 9982).
edge(9982, 9983).
edge(9983, 9984).
edge(9984, 9985).
edge(9985, 9986).
edge(9986, 9987).
edge(9987, 9988).
edge(9988, 9989).
edge(9989, 9990).
edge(9990, 9991).
edge(9991, 9992).
edge(9992, 9993).
edge(9993, 9994).
edge(9994, 9995).
edge(9995, 9996).
edge(9996, 9997).
edge(9997, 9998).
edge(9998, 9999).
edge(9999, 10000).
edge(10000, 0).
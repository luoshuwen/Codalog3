% generate problem of size 1000
reachable(X,Y) :- edge(X,Y).
reachable(X,Y) :- edge(X,Z), reachable(Z,Y).
increasing(X,Y) :- edge(X,Y), lt(X,Y).
increasing(X,Y) :- edge(X,Z), lt(X,Z), increasing(Z,Y).
edge(0, 1).
edge(1, 2).
edge(2, 3).
edge(3, 4).
edge(4, 5).
edge(5, 6).
edge(6, 7).
edge(7, 8).
edge(8, 9).
edge(9, 10).
edge(10, 11).
edge(11, 12).
edge(12, 13).
edge(13, 14).
edge(14, 15).
edge(15, 16).
edge(16, 17).
edge(17, 18).
edge(18, 19).
edge(19, 20).
edge(20, 21).
edge(21, 22).
edge(22, 23).
edge(23, 24).
edge(24, 25).
edge(25, 26).
edge(26, 27).
edge(27, 28).
edge(28, 29).
edge(29, 30).
edge(30, 31).
edge(31, 32).
edge(32, 33).
edge(33, 34).
edge(34, 35).
edge(35, 36).
edge(36, 37).
edge(37, 38).
edge(38, 39).
edge(39, 40).
edge(40, 41).
edge(41, 42).
edge(42, 43).
edge(43, 44).
edge(44, 45).
edge(45, 46).
edge(46, 47).
edge(47, 48).
edge(48, 49).
edge(49, 50).
edge(50, 51).
edge(51, 52).
edge(52, 53).
edge(53, 54).
edge(54, 55).
edge(55, 56).
edge(56, 57).
edge(57, 58).
edge(58, 59).
edge(59, 60).
edge(60, 61).
edge(61, 62).
edge(62, 63).
edge(63, 64).
edge(64, 65).
edge(65, 66).
edge(66, 67).
edge(67, 68).
edge(68, 69).
edge(69, 70).
edge(70, 71).
edge(71, 72).
edge(72, 73).
edge(73, 74).
edge(74, 75).
edge(75, 76).
edge(76, 77).
edge(77, 78).
edge(78, 79).
edge(79, 80).
edge(80, 81).
edge(81, 82).
edge(82, 83).
edge(83, 84).
edge(84, 85).
edge(85, 86).
edge(86, 87).
edge(87, 88).
edge(88, 89).
edge(89, 90).
edge(90, 91).
edge(91, 92).
edge(92, 93).
edge(93, 94).
edge(94, 95).
edge(95, 96).
edge(96, 97).
edge(97, 98).
edge(98, 99).
edge(99, 100).
edge(100, 101).
edge(101, 102).
edge(102, 103).
edge(103, 104).
edge(104, 105).
edge(105, 106).
edge(106, 107).
edge(107, 108).
edge(108, 109).
edge(109, 110).
edge(110, 111).
edge(111, 112).
edge(112, 113).
edge(113, 114).
edge(114, 115).
edge(115, 116).
edge(116, 117).
edge(117, 118).
edge(118, 119).
edge(119, 120).
edge(120, 121).
edge(121, 122).
edge(122, 123).
edge(123, 124).
edge(124, 125).
edge(125, 126).
edge(126, 127).
edge(127, 128).
edge(128, 129).
edge(129, 130).
edge(130, 131).
edge(131, 132).
edge(132, 133).
edge(133, 134).
edge(134, 135).
edge(135, 136).
edge(136, 137).
edge(137, 138).
edge(138, 139).
edge(139, 140).
edge(140, 141).
edge(141, 142).
edge(142, 143).
edge(143, 144).
edge(144, 145).
edge(145, 146).
edge(146, 147).
edge(147, 148).
edge(148, 149).
edge(149, 150).
edge(150, 151).
edge(151, 152).
edge(152, 153).
edge(153, 154).
edge(154, 155).
edge(155, 156).
edge(156, 157).
edge(157, 158).
edge(158, 159).
edge(159, 160).
edge(160, 161).
edge(161, 162).
edge(162, 163).
edge(163, 164).
edge(164, 165).
edge(165, 166).
edge(166, 167).
edge(167, 168).
edge(168, 169).
edge(169, 170).
edge(170, 171).
edge(171, 172).
edge(172, 173).
edge(173, 174).
edge(174, 175).
edge(175, 176).
edge(176, 177).
edge(177, 178).
edge(178, 179).
edge(179, 180).
edge(180, 181).
edge(181, 182).
edge(182, 183).
edge(183, 184).
edge(184, 185).
edge(185, 186).
edge(186, 187).
edge(187, 188).
edge(188, 189).
edge(189, 190).
edge(190, 191).
edge(191, 192).
edge(192, 193).
edge(193, 194).
edge(194, 195).
edge(195, 196).
edge(196, 197).
edge(197, 198).
edge(198, 199).
edge(199, 200).
edge(200, 201).
edge(201, 202).
edge(202, 203).
edge(203, 204).
edge(204, 205).
edge(205, 206).
edge(206, 207).
edge(207, 208).
edge(208, 209).
edge(209, 210).
edge(210, 211).
edge(211, 212).
edge(212, 213).
edge(213, 214).
edge(214, 215).
edge(215, 216).
edge(216, 217).
edge(217, 218).
edge(218, 219).
edge(219, 220).
edge(220, 221).
edge(221, 222).
edge(222, 223).
edge(223, 224).
edge(224, 225).
edge(225, 226).
edge(226, 227).
edge(227, 228).
edge(228, 229).
edge(229, 230).
edge(230, 231).
edge(231, 232).
edge(232, 233).
edge(233, 234).
edge(234, 235).
edge(235, 236).
edge(236, 237).
edge(237, 238).
edge(238, 239).
edge(239, 240).
edge(240, 241).
edge(241, 242).
edge(242, 243).
edge(243, 244).
edge(244, 245).
edge(245, 246).
edge(246, 247).
edge(247, 248).
edge(248, 249).
edge(249, 250).
edge(250, 251).
edge(251, 252).
edge(252, 253).
edge(253, 254).
edge(254, 255).
edge(255, 256).
edge(256, 257).
edge(257, 258).
edge(258, 259).
edge(259, 260).
edge(260, 261).
edge(261, 262).
edge(262, 263).
edge(263, 264).
edge(264, 265).
edge(265, 266).
edge(266, 267).
edge(267, 268).
edge(268, 269).
edge(269, 270).
edge(270, 271).
edge(271, 272).
edge(272, 273).
edge(273, 274).
edge(274, 275).
edge(275, 276).
edge(276, 277).
edge(277, 278).
edge(278, 279).
edge(279, 280).
edge(280, 281).
edge(281, 282).
edge(282, 283).
edge(283, 284).
edge(284, 285).
edge(285, 286).
edge(286, 287).
edge(287, 288).
edge(288, 289).
edge(289, 290).
edge(290, 291).
edge(291, 292).
edge(292, 293).
edge(293, 294).
edge(294, 295).
edge(295, 296).
edge(296, 297).
edge(297, 298).
edge(298, 299).
edge(299, 300).
edge(300, 301).
edge(301, 302).
edge(302, 303).
edge(303, 304).
edge(304, 305).
edge(305, 306).
edge(306, 307).
edge(307, 308).
edge(308, 309).
edge(309, 310).
edge(310, 311).
edge(311, 312).
edge(312, 313).
edge(313, 314).
edge(314, 315).
edge(315, 316).
edge(316, 317).
edge(317, 318).
edge(318, 319).
edge(319, 320).
edge(320, 321).
edge(321, 322).
edge(322, 323).
edge(323, 324).
edge(324, 325).
edge(325, 326).
edge(326, 327).
edge(327, 328).
edge(328, 329).
edge(329, 330).
edge(330, 331).
edge(331, 332).
edge(332, 333).
edge(333, 334).
edge(334, 335).
edge(335, 336).
edge(336, 337).
edge(337, 338).
edge(338, 339).
edge(339, 340).
edge(340, 341).
edge(341, 342).
edge(342, 343).
edge(343, 344).
edge(344, 345).
edge(345, 346).
edge(346, 347).
edge(347, 348).
edge(348, 349).
edge(349, 350).
edge(350, 351).
edge(351, 352).
edge(352, 353).
edge(353, 354).
edge(354, 355).
edge(355, 356).
edge(356, 357).
edge(357, 358).
edge(358, 359).
edge(359, 360).
edge(360, 361).
edge(361, 362).
edge(362, 363).
edge(363, 364).
edge(364, 365).
edge(365, 366).
edge(366, 367).
edge(367, 368).
edge(368, 369).
edge(369, 370).
edge(370, 371).
edge(371, 372).
edge(372, 373).
edge(373, 374).
edge(374, 375).
edge(375, 376).
edge(376, 377).
edge(377, 378).
edge(378, 379).
edge(379, 380).
edge(380, 381).
edge(381, 382).
edge(382, 383).
edge(383, 384).
edge(384, 385).
edge(385, 386).
edge(386, 387).
edge(387, 388).
edge(388, 389).
edge(389, 390).
edge(390, 391).
edge(391, 392).
edge(392, 393).
edge(393, 394).
edge(394, 395).
edge(395, 396).
edge(396, 397).
edge(397, 398).
edge(398, 399).
edge(399, 400).
edge(400, 401).
edge(401, 402).
edge(402, 403).
edge(403, 404).
edge(404, 405).
edge(405, 406).
edge(406, 407).
edge(407, 408).
edge(408, 409).
edge(409, 410).
edge(410, 411).
edge(411, 412).
edge(412, 413).
edge(413, 414).
edge(414, 415).
edge(415, 416).
edge(416, 417).
edge(417, 418).
edge(418, 419).
edge(419, 420).
edge(420, 421).
edge(421, 422).
edge(422, 423).
edge(423, 424).
edge(424, 425).
edge(425, 426).
edge(426, 427).
edge(427, 428).
edge(428, 429).
edge(429, 430).
edge(430, 431).
edge(431, 432).
edge(432, 433).
edge(433, 434).
edge(434, 435).
edge(435, 436).
edge(436, 437).
edge(437, 438).
edge(438, 439).
edge(439, 440).
edge(440, 441).
edge(441, 442).
edge(442, 443).
edge(443, 444).
edge(444, 445).
edge(445, 446).
edge(446, 447).
edge(447, 448).
edge(448, 449).
edge(449, 450).
edge(450, 451).
edge(451, 452).
edge(452, 453).
edge(453, 454).
edge(454, 455).
edge(455, 456).
edge(456, 457).
edge(457, 458).
edge(458, 459).
edge(459, 460).
edge(460, 461).
edge(461, 462).
edge(462, 463).
edge(463, 464).
edge(464, 465).
edge(465, 466).
edge(466, 467).
edge(467, 468).
edge(468, 469).
edge(469, 470).
edge(470, 471).
edge(471, 472).
edge(472, 473).
edge(473, 474).
edge(474, 475).
edge(475, 476).
edge(476, 477).
edge(477, 478).
edge(478, 479).
edge(479, 480).
edge(480, 481).
edge(481, 482).
edge(482, 483).
edge(483, 484).
edge(484, 485).
edge(485, 486).
edge(486, 487).
edge(487, 488).
edge(488, 489).
edge(489, 490).
edge(490, 491).
edge(491, 492).
edge(492, 493).
edge(493, 494).
edge(494, 495).
edge(495, 496).
edge(496, 497).
edge(497, 498).
edge(498, 499).
edge(499, 500).
edge(500, 501).
edge(501, 502).
edge(502, 503).
edge(503, 504).
edge(504, 505).
edge(505, 506).
edge(506, 507).
edge(507, 508).
edge(508, 509).
edge(509, 510).
edge(510, 511).
edge(511, 512).
edge(512, 513).
edge(513, 514).
edge(514, 515).
edge(515, 516).
edge(516, 517).
edge(517, 518).
edge(518, 519).
edge(519, 520).
edge(520, 521).
edge(521, 522).
edge(522, 523).
edge(523, 524).
edge(524, 525).
edge(525, 526).
edge(526, 527).
edge(527, 528).
edge(528, 529).
edge(529, 530).
edge(530, 531).
edge(531, 532).
edge(532, 533).
edge(533, 534).
edge(534, 535).
edge(535, 536).
edge(536, 537).
edge(537, 538).
edge(538, 539).
edge(539, 540).
edge(540, 541).
edge(541, 542).
edge(542, 543).
edge(543, 544).
edge(544, 545).
edge(545, 546).
edge(546, 547).
edge(547, 548).
edge(548, 549).
edge(549, 550).
edge(550, 551).
edge(551, 552).
edge(552, 553).
edge(553, 554).
edge(554, 555).
edge(555, 556).
edge(556, 557).
edge(557, 558).
edge(558, 559).
edge(559, 560).
edge(560, 561).
edge(561, 562).
edge(562, 563).
edge(563, 564).
edge(564, 565).
edge(565, 566).
edge(566, 567).
edge(567, 568).
edge(568, 569).
edge(569, 570).
edge(570, 571).
edge(571, 572).
edge(572, 573).
edge(573, 574).
edge(574, 575).
edge(575, 576).
edge(576, 577).
edge(577, 578).
edge(578, 579).
edge(579, 580).
edge(580, 581).
edge(581, 582).
edge(582, 583).
edge(583, 584).
edge(584, 585).
edge(585, 586).
edge(586, 587).
edge(587, 588).
edge(588, 589).
edge(589, 590).
edge(590, 591).
edge(591, 592).
edge(592, 593).
edge(593, 594).
edge(594, 595).
edge(595, 596).
edge(596, 597).
edge(597, 598).
edge(598, 599).
edge(599, 600).
edge(600, 601).
edge(601, 602).
edge(602, 603).
edge(603, 604).
edge(604, 605).
edge(605, 606).
edge(606, 607).
edge(607, 608).
edge(608, 609).
edge(609, 610).
edge(610, 611).
edge(611, 612).
edge(612, 613).
edge(613, 614).
edge(614, 615).
edge(615, 616).
edge(616, 617).
edge(617, 618).
edge(618, 619).
edge(619, 620).
edge(620, 621).
edge(621, 622).
edge(622, 623).
edge(623, 624).
edge(624, 625).
edge(625, 626).
edge(626, 627).
edge(627, 628).
edge(628, 629).
edge(629, 630).
edge(630, 631).
edge(631, 632).
edge(632, 633).
edge(633, 634).
edge(634, 635).
edge(635, 636).
edge(636, 637).
edge(637, 638).
edge(638, 639).
edge(639, 640).
edge(640, 641).
edge(641, 642).
edge(642, 643).
edge(643, 644).
edge(644, 645).
edge(645, 646).
edge(646, 647).
edge(647, 648).
edge(648, 649).
edge(649, 650).
edge(650, 651).
edge(651, 652).
edge(652, 653).
edge(653, 654).
edge(654, 655).
edge(655, 656).
edge(656, 657).
edge(657, 658).
edge(658, 659).
edge(659, 660).
edge(660, 661).
edge(661, 662).
edge(662, 663).
edge(663, 664).
edge(664, 665).
edge(665, 666).
edge(666, 667).
edge(667, 668).
edge(668, 669).
edge(669, 670).
edge(670, 671).
edge(671, 672).
edge(672, 673).
edge(673, 674).
edge(674, 675).
edge(675, 676).
edge(676, 677).
edge(677, 678).
edge(678, 679).
edge(679, 680).
edge(680, 681).
edge(681, 682).
edge(682, 683).
edge(683, 684).
edge(684, 685).
edge(685, 686).
edge(686, 687).
edge(687, 688).
edge(688, 689).
edge(689, 690).
edge(690, 691).
edge(691, 692).
edge(692, 693).
edge(693, 694).
edge(694, 695).
edge(695, 696).
edge(696, 697).
edge(697, 698).
edge(698, 699).
edge(699, 700).
edge(700, 701).
edge(701, 702).
edge(702, 703).
edge(703, 704).
edge(704, 705).
edge(705, 706).
edge(706, 707).
edge(707, 708).
edge(708, 709).
edge(709, 710).
edge(710, 711).
edge(711, 712).
edge(712, 713).
edge(713, 714).
edge(714, 715).
edge(715, 716).
edge(716, 717).
edge(717, 718).
edge(718, 719).
edge(719, 720).
edge(720, 721).
edge(721, 722).
edge(722, 723).
edge(723, 724).
edge(724, 725).
edge(725, 726).
edge(726, 727).
edge(727, 728).
edge(728, 729).
edge(729, 730).
edge(730, 731).
edge(731, 732).
edge(732, 733).
edge(733, 734).
edge(734, 735).
edge(735, 736).
edge(736, 737).
edge(737, 738).
edge(738, 739).
edge(739, 740).
edge(740, 741).
edge(741, 742).
edge(742, 743).
edge(743, 744).
edge(744, 745).
edge(745, 746).
edge(746, 747).
edge(747, 748).
edge(748, 749).
edge(749, 750).
edge(750, 751).
edge(751, 752).
edge(752, 753).
edge(753, 754).
edge(754, 755).
edge(755, 756).
edge(756, 757).
edge(757, 758).
edge(758, 759).
edge(759, 760).
edge(760, 761).
edge(761, 762).
edge(762, 763).
edge(763, 764).
edge(764, 765).
edge(765, 766).
edge(766, 767).
edge(767, 768).
edge(768, 769).
edge(769, 770).
edge(770, 771).
edge(771, 772).
edge(772, 773).
edge(773, 774).
edge(774, 775).
edge(775, 776).
edge(776, 777).
edge(777, 778).
edge(778, 779).
edge(779, 780).
edge(780, 781).
edge(781, 782).
edge(782, 783).
edge(783, 784).
edge(784, 785).
edge(785, 786).
edge(786, 787).
edge(787, 788).
edge(788, 789).
edge(789, 790).
edge(790, 791).
edge(791, 792).
edge(792, 793).
edge(793, 794).
edge(794, 795).
edge(795, 796).
edge(796, 797).
edge(797, 798).
edge(798, 799).
edge(799, 800).
edge(800, 801).
edge(801, 802).
edge(802, 803).
edge(803, 804).
edge(804, 805).
edge(805, 806).
edge(806, 807).
edge(807, 808).
edge(808, 809).
edge(809, 810).
edge(810, 811).
edge(811, 812).
edge(812, 813).
edge(813, 814).
edge(814, 815).
edge(815, 816).
edge(816, 817).
edge(817, 818).
edge(818, 819).
edge(819, 820).
edge(820, 821).
edge(821, 822).
edge(822, 823).
edge(823, 824).
edge(824, 825).
edge(825, 826).
edge(826, 827).
edge(827, 828).
edge(828, 829).
edge(829, 830).
edge(830, 831).
edge(831, 832).
edge(832, 833).
edge(833, 834).
edge(834, 835).
edge(835, 836).
edge(836, 837).
edge(837, 838).
edge(838, 839).
edge(839, 840).
edge(840, 841).
edge(841, 842).
edge(842, 843).
edge(843, 844).
edge(844, 845).
edge(845, 846).
edge(846, 847).
edge(847, 848).
edge(848, 849).
edge(849, 850).
edge(850, 851).
edge(851, 852).
edge(852, 853).
edge(853, 854).
edge(854, 855).
edge(855, 856).
edge(856, 857).
edge(857, 858).
edge(858, 859).
edge(859, 860).
edge(860, 861).
edge(861, 862).
edge(862, 863).
edge(863, 864).
edge(864, 865).
edge(865, 866).
edge(866, 867).
edge(867, 868).
edge(868, 869).
edge(869, 870).
edge(870, 871).
edge(871, 872).
edge(872, 873).
edge(873, 874).
edge(874, 875).
edge(875, 876).
edge(876, 877).
edge(877, 878).
edge(878, 879).
edge(879, 880).
edge(880, 881).
edge(881, 882).
edge(882, 883).
edge(883, 884).
edge(884, 885).
edge(885, 886).
edge(886, 887).
edge(887, 888).
edge(888, 889).
edge(889, 890).
edge(890, 891).
edge(891, 892).
edge(892, 893).
edge(893, 894).
edge(894, 895).
edge(895, 896).
edge(896, 897).
edge(897, 898).
edge(898, 899).
edge(899, 900).
edge(900, 901).
edge(901, 902).
edge(902, 903).
edge(903, 904).
edge(904, 905).
edge(905, 906).
edge(906, 907).
edge(907, 908).
edge(908, 909).
edge(909, 910).
edge(910, 911).
edge(911, 912).
edge(912, 913).
edge(913, 914).
edge(914, 915).
edge(915, 916).
edge(916, 917).
edge(917, 918).
edge(918, 919).
edge(919, 920).
edge(920, 921).
edge(921, 922).
edge(922, 923).
edge(923, 924).
edge(924, 925).
edge(925, 926).
edge(926, 927).
edge(927, 928).
edge(928, 929).
edge(929, 930).
edge(930, 931).
edge(931, 932).
edge(932, 933).
edge(933, 934).
edge(934, 935).
edge(935, 936).
edge(936, 937).
edge(937, 938).
edge(938, 939).
edge(939, 940).
edge(940, 941).
edge(941, 942).
edge(942, 943).
edge(943, 944).
edge(944, 945).
edge(945, 946).
edge(946, 947).
edge(947, 948).
edge(948, 949).
edge(949, 950).
edge(950, 951).
edge(951, 952).
edge(952, 953).
edge(953, 954).
edge(954, 955).
edge(955, 956).
edge(956, 957).
edge(957, 958).
edge(958, 959).
edge(959, 960).
edge(960, 961).
edge(961, 962).
edge(962, 963).
edge(963, 964).
edge(964, 965).
edge(965, 966).
edge(966, 967).
edge(967, 968).
edge(968, 969).
edge(969, 970).
edge(970, 971).
edge(971, 972).
edge(972, 973).
edge(973, 974).
edge(974, 975).
edge(975, 976).
edge(976, 977).
edge(977, 978).
edge(978, 979).
edge(979, 980).
edge(980, 981).
edge(981, 982).
edge(982, 983).
edge(983, 984).
edge(984, 985).
edge(985, 986).
edge(986, 987).
edge(987, 988).
edge(988, 989).
edge(989, 990).
edge(990, 991).
edge(991, 992).
edge(992, 993).
edge(993, 994).
edge(994, 995).
edge(995, 996).
edge(996, 997).
edge(997, 998).
edge(998, 999).
edge(999, 1000).
edge(1000, 0).
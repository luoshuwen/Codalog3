% generate problem of size 10
reachable(X,Y) :- edge(X,Y,Z).
reachable(X,Y) :- edge(X,Z), reachable(Z,Y).
same_clique(X,Y) :- reachable(X,Y), reachable(Y,X).
%edge(X,Y):-edge(X,Y).
edge(0, 1).
edge(1, 2).
edge(2, 'A b').
edge('A b',0).
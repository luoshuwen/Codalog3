%P.cdl
p(X,N):-p(X,Z),p(Z,Y).
p(X,Y):-e(X,Y).%,X>1.
e(1,2).
e(2,X). 
%e(3,1).